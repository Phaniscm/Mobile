63e4144b
31c30494
700f7e72
31c3300c
2000341c
313c68d2
63e4138b
31c30494
700f7e92
31c3300c
211c4006
32834000
10546007
0540503c
363c31c3
7072145b
3bc3700f
13546007
108c353c
786e69c3
503c01d3
31c30340
139b363c
700f6d72
05d20bc3
108c353c
644e19c3
32c3500c
611cc006
36034000
0f8b133c
313c32c3
700f0f9b
01d36006
024f073c
2b9d013c
0034323c
02946067
4025e205
f5944207
1d810133
608515e1
fc946407
40060073
0026fd93
0f56f076
00000804
50c37016
d1e9848c
1771005c
7fe530c3
0b3563e4
301c0116
311c0b84
6c0c0000
00b1001c
80563664
0cc7363c
0584255c
708b2d00
110b65ee
512b054f
44cc450f
23837f86
10c944cf
341c30c3
32a30003
50cb64cf
1586255c
44ee514b
65d26409
03546047
13c6255c
0e560006
00000804
fe96f016
1233705c
59e9c48c
17c7323c
0564205c
79c92d00
00f4433c
094b233c
090b333c
34546007
24944007
023c4026
0077400d
07a9315c
007703a3
00210f5c
07ad015c
0080343c
300d323c
32a347ec
343c67ef
658000c7
035c188b
133c07e6
58ab1000
336432c3
02356407
442e4406
215c04b3
40070ba3
60262194
315c3423
622c0ba6
39e96c2c
3664588b
4ef202f3
34236026
403723e3
07a9315c
40372383
00010f5c
07ad015c
60260133
33e33423
0ba3215c
315c3283
37c40ba6
f88c033c
0f560296
00000804
ff96f016
e06c50c3
625c448c
28eb0034
341c31c3
64f2000f
780e68ab
20860373
9fcc2037
43e62026
46646006
355c20c3
606517c4
31833f86
61806205
2c0e2006
2c0e380b
2c2e2006
0404375c
12c305c3
00063664
0f560196
00000804
ff963016
29e2648c
320b413c
0b04301c
0000311c
523c4c09
a0370010
00010f5c
47f20c0d
311c6386
4c0f2010
4c0f6085
0034013c
1b540027
004706d2
00672e54
06733b94
09b483e7
211c4386
280c2010
34236026
02b331a3
211c4406
080c2010
01f4143c
31236026
017330a3
0cb483e7
211c4386
280c2010
400d303c
318333e3
480c680f
44060333
2010211c
343c280c
303c01f4
fe73300d
311c6386
a0062010
6085ac0f
0113ac0f
311c6386
1fe62010
60850c0f
00060c0f
0c560196
00000804
648c7016
880c40ec
52c34d09
123c4d29
ad4942ac
ad6965c3
432c253c
00064664
08040e56
1f36f016
70c3ff96
c48ca1c3
0011865c
60ac2070
a2ac4c4c
0021b65c
c23c38c3
4bc33a1d
04c4355c
c6645180
78cb0ad2
80378006
89ec29c3
202607c3
466428c3
724c49c3
1a3c07c3
36640040
f8760196
08040f56
0aa3105c
105c31c3
31a30ac3
0ab3105c
305c31a3
08040a96
1f36f016
70c3ff96
4010c2c3
6cd03ac3
cc4c60ac
9549a48c
341c34c3
946c0001
343c6ad2
64d20c8b
07c4365c
365c0173
011307a4
240b443c
0044343c
365c65d2
36640784
855c0433
d5290041
0034943c
0014343c
60cc64d2
36646dcc
211c4006
40378000
8c8c3bc3
2cc30ac3
28c33500
466436c3
0024393c
66d20026
706c4bc3
36641c0c
01960026
0f56f876
00000804
50c3f016
72c341c3
6dcc60cc
908c3664
cfec746c
338005c3
71295109
540c6664
6c6c68cc
366402c3
0f560006
00000804
0336f016
60c3ff96
0070a0ac
70eb848c
941c93c3
39c30004
744c66f2
07e4335c
07133664
928494c3
573cf109
a037080c
8fcc38c3
40662026
46646006
365c10c3
531c17c4
093500ff
5f866065
61803283
40724ceb
ac4e4cee
17c4365c
9f866065
62053483
40060580
343c49c3
6112259d
8000401c
2010411c
8c0b6e00
271d403c
27e44025
48c3f214
0404345c
366406c3
01960006
0f56c076
00000804
0136f016
82c350c3
cccc600c
50eb848c
341c32c3
733c000f
341c0034
67d20001
0a83305c
60cc64f2
36646dcc
0424365c
28c31109
40063100
373c3664
64d20024
140c786c
00263664
0f568076
00000804
ff96f016
72c340c3
648cc06c
24066c49
bbcc2037
23c32026
56646006
345c20c3
606517c4
31833f86
61807d80
27a3145c
145c2c0e
2c2e27b3
0404365c
12c304c3
00063664
0f560196
00000804
3f36f016
80c3fd96
006c32c3
448c00b7
0051c25c
28ebc909
541c51c3
a0770003
0002c31c
69800e94
b35cec0b
a35c0013
433c0023
563c0060
901c0067
02730000
0001c31c
a0060854
b5c375c3
95c3a5c3
013345c3
100c563c
0063925c
b7c3e006
47c3a7c3
4097a037
08c3abd0
42862026
d6646006
08c3d0c3
17c4305c
00ff531c
60650a35
32835f86
61800dc3
40724ceb
ac4e4cee
315c18c3
606517c4
32835f86
0dc36205
2057a180
341c31c3
66d20001
68cc28c3
08c36dcc
c31c3664
21940002
080c373c
8000101c
2010111c
3b3c0c80
2c80080c
080c3a3c
8000201c
2010211c
25c36d00
b00b0193
b04ba00e
a40bac0e
ac0ba82e
40c5a84e
dfe580c5
0473d5f2
c31c15c3
1f940001
29c30393
1800221c
100c323c
8000501c
2010511c
6c0b6e80
323c640e
001c100c
011c8002
6c002010
642e6c0b
dfe52085
0010393c
936493c3
e494c007
35c3a057
0002341c
08c367d2
4ccc600c
03c3486c
20972664
0404315c
1dc308c3
00063664
fc760396
08040f56
3f36f016
d0c3ff96
648ca0ac
843c8c6c
683c240b
c6d20044
335c744c
36640764
143c13b3
2037250b
0051b35c
0041c35c
b31c4d00
0a940002
a25ce80b
925c0013
423c0023
56c30060
b31c01f3
07540001
76c356c3
96c3a6c3
00d346c3
42c3accb
a6c376c3
683c96c3
383c0034
66d20014
64cc1dc3
0dc36dcc
700b3664
ffff201c
0000211c
30e402c3
20171a94
341c31c3
60070001
502b1394
62c64ad2
4105311c
23644c0b
0018251c
01134c0e
211c42c6
680b4105
fff7341c
8085680e
0002b31c
373c1d94
501c080c
511c8000
0e802010
080c3a3c
393c2e80
4e80080c
700b0193
b02b600e
704ba40e
80c5680e
fff03c3c
c364c3c3
74f23cc3
b31c04d3
23940001
201c03f3
35001800
100c313c
8000001c
2010011c
700b4c00
313c680e
101c100c
111c8002
4c802010
680e702b
3c3c8085
c3c3ffe0
353cc364
53c30010
3cc35364
e0946007
0024363c
68d20026
740c5dc3
486c4ccc
266403c3
01960026
0f56fc76
00000804
ff96f016
605c50c3
800c0544
0909448c
0624145c
0229315c
03546027
04946127
60376006
48c90073
7f5c4037
e6ed0001
303c79ac
79af20db
05b40027
745ce026
009303d5
345c6046
104c03d5
2cbc16c3
00070880
74cc1294
05c36dcc
765c3664
27c301c1
0001241c
201c43d2
70cc4000
04c36d8c
366416c3
01960026
08040f56
0136f016
705c40c3
c06c0544
0270a00c
17c3144c
08802cbc
01160ad2
0b84301c
0000311c
0c666c0c
80563664
0444365c
366404c3
6c0c74ec
17c305c3
365c3664
04c304e4
365c3664
04c304a4
365c3664
04c304c4
28c33664
04c3686c
00063664
0f568076
00000804
305c20c3
105c0ae4
31830b04
125c03c3
01830b24
1341125c
087374bc
00000804
105c31e3
31830b24
0b27305c
0904aabc
00000804
0b24305c
305c31a3
aabc0b27
08040904
0b27105c
0904aabc
00000804
105c31e3
31830b04
0b07305c
0904aabc
00000804
0b04305c
305c31a3
aabc0b07
08040904
0b07105c
0904aabc
00000804
105c31e3
31830ae4
0ae7305c
0904aabc
00000804
0ae7105c
0904aabc
00000804
800c1016
0d09648c
40074cc9
345c1694
66d20d91
311c6506
4c0e4020
658600d3
4140311c
4c0f4086
08959cbc
345c0004
60070d91
03932254
0e944027
0d91245c
311c6586
40074140
65061b54
4020311c
4c0e4006
406702f3
301c0894
311c0448
4c0c2010
01b34072
0d91245c
650646d2
4020311c
fdd34206
311c6606
40864140
70cc4c0f
045c6d4c
36640624
08560006
00000804
40c33016
a4c9248c
2394a007
021c62ac
22050234
05a4235c
08cbb0bc
11a3345c
345c6bd2
345c0a01
545c12c5
62460a07
0447345c
006602b3
0fe4301c
0000311c
b4bc2cac
345c0873
345c12c1
01130a07
305c6086
606c0a6d
05e4335c
00063664
08040c56
0424205c
11544007
04e4325c
325c6f72
600604e7
04c6325c
301c0066
311c0fe4
2cac0000
0873b4bc
00000804
40c33016
ad09648c
035c600c
09d20361
301c0066
311c0fe4
2cac0000
0873b4bc
5694a007
145c2026
301c0a86
311c8606
0c0b2010
241c20c3
2364effd
4c0e4072
8604201c
2010211c
31c3280b
1003351c
201c680e
211c8004
680b2010
680e6d72
0620221c
30c3080b
feff341c
201c680e
211c8622
280b2010
341c31c3
680eff8f
82c2201c
2010211c
6072680b
101c680e
111c8644
440b2010
341c32c3
3364fffb
640e6072
8642301c
2010311c
0c0e0206
860c201c
2010211c
30c3080b
0007351c
440b680e
351c32c3
640e0005
a02708b3
00064354
0a86045c
8604201c
2010211c
31c3280b
effc341c
4045680e
30c3080b
effc341c
201c680e
211c8004
280b2010
341c31c3
680edfff
0620221c
6872680b
201c680e
211c8622
080b2010
351c30c3
680e0070
82c2201c
2010211c
31c3280b
fffe341c
221c680e
080b0382
341c30c3
680efffa
860c201c
2010211c
31c3280b
0007351c
0026680e
08040c56
40c31016
2d09648c
2d2921c3
412c313c
0c76305c
0010341c
8ebc65d2
045c0895
002615a7
08040856
0136f016
70c3f996
19e9c48c
303c0177
275c0cc7
ad000584
0641355c
0d946027
602778a9
01160a94
0b84301c
0000311c
07666c0c
80563664
21b738a9
06942027
00c13f5c
0645355c
81970a13
004704c3
155c3f94
20070641
0014a2dc
63d27409
14946047
1504375c
04c38c09
01371fe5
00811f5c
375c2c0d
2c091504
275c27f2
686c0604
095b313c
7409686f
0a946067
14e1375c
9fe543c3
0f5c80f7
075c0061
7eac14e5
135c05c3
9cbc0464
375c08cb
2c091504
200720b7
0011a4dc
00412f5c
375c4d0d
4f5c1504
8c2d0041
01972213
206710c3
01160a54
0b84301c
0000311c
07e66c0c
80563664
32c358eb
000f341c
00c7333c
04e4475c
742f6e00
140d1909
342d3929
548e590b
74ae792b
94ce994b
14ee196b
350e398b
552e59ab
754e79cb
94cf990c
15ce1a4b
35ee3a6b
550f594c
752f796c
954f998c
16ce1b6b
135c7c0c
25f20361
275c5b8b
00931586
375c6286
74091586
604766d2
14eb0454
13c6075c
748b54ab
813c2157
2067180c
223c19b4
608681ac
2010311c
34cb4c0f
2c0f6085
011c0186
400c2010
00ff301c
33e33823
213c3283
2823408c
600f32a3
223c0353
620681ac
2010311c
14cb4c0f
0c0f6085
411c8306
500c2010
fe00183c
00ff301c
33e33123
203c3283
2123408c
700f32a3
60277409
60670354
2f5c0c94
275c00a1
7b4b147d
375c6a12
865c12e7
00f301a3
175c1b4b
5cbc1771
80c30a7c
1504375c
85d28c09
63d27409
14946047
08c4301c
2010311c
483c0c11
7dcc500c
07c36c0c
402614c3
50203664
08c8301c
2010311c
74094c0f
604763d2
375c4e94
40261504
375c4d0d
9b4b1504
375c8c2e
0f5c1504
0d4d00a1
602778a9
375c0a94
4c091504
802542c3
0f5c8077
0c0d0021
000d831c
301c0e35
311c08e0
201c2010
4c0f2ee0
1504375c
1f40401c
04b38c2f
ff90383c
0b84001c
0000011c
17b460a7
3e87183c
c180213c
08e0301c
2010311c
275c4c0f
401c1504
6600ec78
0116682f
001c600c
366400a4
00f38056
600c0116
00a4001c
80563664
60677409
175c0a94
21c314e1
40374025
00013f5c
14e5375c
07960006
0f568076
00000804
40c3f016
0524505c
0504305c
63c3740f
000613c3
0200201c
6006440e
345c642e
606517c4
3783ff86
e006442c
0025ed61
345c2105
03e40941
f42fee14
6dcc70cc
366404c3
311c6a86
ffe62010
72acec0f
2d8c05c3
08cb9cbc
0113a006
06c3a025
0424125c
08cb9cbc
345cc105
52ac0941
f51453e4
0e00043c
04e4125c
08cb9cbc
211c4006
680c2010
dffe701c
680f3783
0400221c
6092680c
301c680f
311c0fe4
6d8c0000
0b30001c
0000011c
301c3664
311c0246
20062020
0f562c0e
00000804
0336f016
905c50c3
e48c0664
31c33ca9
0003341c
6cf25cab
205c32e3
32830ac3
0ac6305c
31a33c8b
0ac6305c
32e30173
0ab3205c
305c3283
3c8b0ab6
305c31a3
746c0ab6
05c36e8c
5ceb3664
0b46255c
83c37ceb
83a37cab
383cc006
341c608d
6dd20001
0070463c
155c04c3
00bc1341
04c30873
1341155c
0872a2bc
c107c025
7cc9ed94
0ad6355c
323c5cc9
60070014
19c31254
341c640c
6dd20001
0024323c
1341155c
028665d2
0872d0bc
02860093
087300bc
c0760006
08040f56
0136f016
60c3ff96
62ac0070
05c4335c
0440533c
18c3a037
212687cc
60064466
70c34664
17c4365c
5f866065
5aac3283
04a4125c
81806c80
15c304c3
08cb9cbc
1384365c
0a24235c
365c500f
535c1384
b04e09c3
1384365c
306e2fcb
200606c3
08e73abc
06c3108e
3abc2026
10ae08e7
204606c3
08e73abc
106f0364
0b1c301c
0000311c
508f4c0c
0b08301c
0000311c
b0afac0c
0448301c
2010311c
70cf6c0c
008c301c
2010311c
70ef6c0c
790c201c
2010211c
710f680c
712f680c
714f680c
335c780c
2e0c0624
04c3316f
400614c3
06a4365c
accb6d00
4785a70e
231c2045
f79402d0
365c4006
6d0006a4
a24fac8c
06a4365c
2cec6d00
4785226f
231c0105
f29402d0
2524365c
545cacec
165c0547
145c0a93
265c0566
245c0ab3
365c0576
345c0ac3
565c0586
545c0aa3
7aac0596
05c4335c
31833f86
04c39180
0644165c
b0bc4086
043c08cb
101c0040
111c0dbc
48060000
08cbb0bc
325c28c3
06c30404
366417c3
80760196
08040f56
0bb4301c
0000311c
335c6c0c
0ccc1804
00000804
0336f016
60c3fc96
72c301c3
a48c83c3
17a4165c
235c7aac
74a904c4
95e960b7
3f5c80f7
305c0061
7dac01ed
0eb460e7
343c80d7
465c17c7
6e000564
341c6c0c
60070002
000ad4dc
74ca00b3
83dc6007
946b000a
341c34c3
64d20010
6f72620c
94cb620f
341c34c3
64d24000
7672620c
94cb620f
341c34c3
64d21000
7e72620c
6006620f
27c5365c
34c3946b
0040341c
602664d2
27c5365c
34c39449
0001341c
10946007
609761af
806543c3
43837f86
4f5c8077
405c0021
3f5c01dd
305c0041
800601e5
946b818f
341c34c3
80860001
744c6fd2
7609622f
0246305c
0a61465c
762986d2
0824401c
02546067
746b8486
941c93c3
39c30200
817262d2
93c37469
0010941c
67d239c3
6c806100
105c2c29
00b301fd
0a01265c
01fd205c
32c3546b
60073164
323c2415
60078004
87721f54
341c32c3
746efffb
4004323c
9d7262d2
0544365c
265c6dac
133c04e4
6829424b
0c5413e4
25c1365c
921c93c3
9f5c0001
1f5c0007
165c0001
887225c5
61277dac
620c0494
620f7172
323c546b
62d20044
323c8372
62d20024
54699272
0204323c
997262d2
0404323c
987267d2
620c00b3
620f6472
620ceaf3
620f34a3
604e6006
604c606e
00ff401c
9fff411c
7f923483
34cb604f
0266105c
00412f5c
18c3410d
7aac1364
235c838b
71200484
604c4ca0
6c1b323c
7aac604f
235c80cb
71200484
60ce6ca0
48c37aac
0484135c
408c7080
608f6d00
c0760496
08040f56
42321016
46d26006
85e18181
60855fe5
0856ff73
00000804
41321016
080c323c
01802580
7fc56006
85e245d2
5fe581c1
0856ff73
00000804
40c31016
11cb213c
08544027
104b013c
00064ed2
0b944047
313c00d3
033c0074
00b30040
07f4313c
00c0033c
335c700c
604703d1
1f850294
08040856
0136f016
51c340c3
115c72c3
313c0279
205c0cc7
cd000584
323c560c
63d20204
0a33362c
341c78cc
63d20001
0973394c
0024323c
01166ad2
0b84301c
0000311c
02e66c0c
80563664
01e9155c
17c7313c
0564145c
025c4c80
760c0463
111c2006
31834000
125c6fd2
31c307a9
01f1155c
341c3143
66d20001
0443125c
033c6080
101c0010
325c008b
65d20403
0520303c
359d123c
5804313c
331c182c
04540100
6c32604b
004b01d3
325c0ed2
602702a9
60060694
0006311c
00b313a3
608c303c
80ac133c
5804313c
331c64d2
09940080
0a61245c
782c46f2
6c326c4b
241b133c
613c362f
cef25804
0ca3245c
341c32c3
68d20001
201c31c3
211c0200
32a30010
700c762f
0624335c
40074e09
722c3754
04c36ccc
20c33664
fff0363c
033c7f32
323c380c
64120330
640b3180
0246355c
200c323c
633c7180
78683340
27a6345c
245c440b
345c27b6
600727e1
245c1794
400727d1
201c1394
211c3a01
7d001008
442b6112
0c0e02a3
3a68101c
1008111c
233c7c80
780b080c
355c680e
6bf20243
00d2201c
0246255c
27a6345c
0243355c
27b6345c
0f568076
00000804
40c37016
62c351c3
422c6364
13c348cc
145c2664
200727e1
303c1654
7180200c
19a3135c
241c21c3
303c0007
64120330
6c2b7180
323c6c12
263c49ac
32a31ff4
03d3742f
27d1245c
1a544007
303c15c3
1180200c
19b1605c
341c36c3
605c001f
263c19c3
213c29ac
345c027e
68d227d9
19e4305c
812c233c
7032440f
0e56744f
00000804
3f36f016
b0c3f796
259081c3
460ca630
2004323c
09c36bd2
0623a05c
0633505c
0800601c
0010611c
19c301b3
04f3015c
341c30c3
a33c1fff
c0060040
0010611c
18c3a026
0243115c
323c21b7
6dd20024
025c28c3
20c30279
0cc7323c
005c0bc3
8c000584
01934006
215c18c3
12c301e9
17c7313c
005c0bc3
4c000564
cd3c8a8c
3c3c5804
7fe51806
f88c733c
c31ce4f2
07940400
0594a027
09c32286
009322ce
39c30086
38c30ece
313c2e0c
61370024
31c36ef2
011c0006
30830040
67f260f7
2004313c
d17263d2
d0720053
a027e7d2
36c30594
63c37192
313cd072
60070104
01174f54
15540007
05c4245c
200632c3
4000111c
333c3103
133c0f8b
023c280c
343c2a0b
6c800340
29c36232
01936b0e
044f123c
7f3231e3
013c6512
6980288b
19c36232
cc72670e
0014303c
353c66d2
2ac3180c
02f36980
0104303c
651c68d2
353ca000
1ac3200c
01b36580
00a4303c
08c36cd2
01f9305c
02b46027
cf72de72
00c03a3c
0173a3c3
0044303c
00401a3c
651c64d2
00536000
a1c3ce72
28c3a364
313c2a0c
62d20084
313cd672
62d21004
6206dd72
0cc361f7
414603f2
2d3c41f7
c2c3808c
31c3c364
011c0006
30830400
c27262d2
18043d3c
0fff241c
392c333c
644f19c3
225c2bc3
45f227e1
335c3bc3
6bd227d1
622c0bc3
193c8f2c
61970080
3dc323c3
00b34664
68126197
606f09c3
115c1bc3
25d227e1
68126197
688f29c3
7ff45d3c
620c08c3
0002341c
d7c3e006
15946007
662c1bc3
36c38cec
211c4006
32830001
62f221c6
05c32306
3f3c2cc3
46640220
61d70364
d7c3e180
a1775364
622c0bc3
05c38cec
2cc31ac3
02203f3c
28c34664
0256025c
32c34a0c
011c0006
30830008
b49256c3
18946007
341c32c3
66d22000
737236c3
b69253c3
19c301f3
56c3e66e
28c3b572
341c6a0c
66d20001
600656c3
08a0311c
08c353a3
2006620c
0020111c
68d23183
005c2dc3
68000253
315c18c3
2bc30286
cf5c6a2c
0f5c0006
0f5c0113
20060026
8f4c20b7
0180093c
12c34157
35c32ac3
38c34664
32c34e0c
011c0006
30830002
551c63d2
323c0042
6ad20804
32c3a772
111c2006
31832000
551c63d2
28c300c2
01f9325c
02b46027
19c3be72
0996a54f
0f56fc76
00000804
3f36f016
70c3f996
40f7c1c3
115c43c3
213701e9
0564b05c
125c2cc3
21c30279
0cc7323c
105cd3c3
d1840584
2f5c4006
3cc300d6
1dc3cd8c
6c4b642c
533c6c32
452c800c
600c52a3
0624335c
20072e09
4d894e54
4b944007
6ccc622c
366415c3
5804353c
7f327fe5
380c933c
0330303c
3d806412
0003815c
27e1375c
24946007
27d1275c
20944007
3a01201c
1008211c
a33c7100
2ac3080c
3364680b
333c442b
39a3412c
1ac33364
201c640e
211c3a74
71001008
080c233c
200c303c
335c7d80
680e19a3
101c02f3
111c3a01
70801008
080c133c
2364440b
0330303c
7d806412
323c0c2b
3364402c
0093640e
815c1cc3
353c0243
a3c3808c
253ca364
341c1804
323c0fff
79cf39ac
27d1375c
075c64f2
0ad227e1
8f2c7e2c
163c07c3
28c30380
466435c3
383c0093
79ef400c
27e1175c
383c24d2
7a0f400c
7ff4953c
5804353c
41774206
614663f2
00d76177
202710c3
41172b94
17c7323c
61800bc3
00b4101c
02c6165c
0243235c
02e6265c
0253035c
02f6065c
0263135c
0306165c
8cec7e2c
21c609c3
3f3c2ac3
466401a0
b364b0c3
4000301c
02a6365c
065c0206
801c02b6
62860005
101c0233
165c00c4
201c02c6
265c8000
614602a6
02b6365c
0002801c
b01c61c6
59c30000
93c35364
7e2c9364
05c38cec
2ac319c3
01a03f3c
7e2c4664
0006af5c
00d31f5c
00261f5c
40b74006
063c8f4c
15c30480
600629c3
21574664
005c0cc3
64000253
365c3b84
383c02d6
1dc302c0
163c248b
383c371d
2dc302d0
263c48ab
383c371d
0dc302e0
063c00cb
0796371d
0f56fc76
00000804
7d72602c
602f6f92
602e6006
622b600e
620b69f2
616b6af2
614b6bf2
60ab6cf2
620b6df2
620e6e72
6e72616b
614b616e
614e6e72
6e7260ab
608b60ae
608e6e72
00000804
40c37016
682c03c3
aa0b602f
c96ba22e
694bc20e
a8ab616e
c88ba14e
01e1515c
60ae7aa0
01d9315c
c92c608e
68ecc14f
a8cc612f
c88ca0ef
315cc0cf
a86c01e1
608f6e80
c006660c
1000611c
64d23683
606f65ac
a86c0073
722ca06f
36646d0c
08040e56
105cfe96
21c30159
40375fe5
00011f5c
2f5c2077
205c0021
618c015d
1a1d033c
08040296
0159205c
0b0d323c
7f327fe5
080403c3
ff967016
62c340c3
acec622c
230601c3
3f3c4006
56640020
536450c3
1771245c
1504145c
68000549
323c8f20
4383fff0
0a12042b
5cbc12c3
343c0a7c
1580028d
0e560196
00000804
fe967016
61c340c3
0544305c
4dac20cc
424b323c
244b223c
00062f5c
40774006
20a6a5ec
56644026
201c722c
211c2a18
4d2f0012
6d2c722c
16c304c3
02963664
08040e56
ff961016
205c40c3
616c0149
2b9d133c
0149205c
602532c3
2f5c6037
205c0001
2af2014d
301c0116
311c0b84
6c0c0000
366404e6
245c8056
345c0149
23e40141
01160a35
0b84301c
0000311c
05066c0c
80563664
08560196
00000804
ff963016
51c340c3
0159205c
240c618c
2b9d133c
0159205c
602532c3
1f5c6037
105c0001
740c015d
01166af2
0b84301c
0000311c
05266c0c
80563664
540f4006
0159245c
0151345c
0a3523e4
301c0116
311c0b84
6c0c0000
36640546
01968056
08040c56
ff967016
52c341c3
245c238c
323c0279
605c0cc7
6f000584
345c4c09
6bd201f9
0a61605c
633cc8f2
c037fff0
00010f5c
01fd045c
1494a007
8006720c
0840411c
c0063483
0800611c
30e406c3
40272694
40670354
648c2294
648f6025
c48b03d3
602536c3
045c648e
000701f9
442b1694
602532c3
64cb642e
03546027
cbf2c46b
30c3046b
23c36025
446e2364
32e4644b
444e0234
c4cec026
0e560196
00000804
fe967016
41c360c3
536452c3
01e9315c
660c6077
660f6072
6dcc622c
366425c3
32c3520c
111c2006
31830800
15546007
01f9345c
a2d263f2
323ca046
60370204
7a8c6cf2
06c38c0c
5f5c15c3
25c30021
00015f5c
466435c3
0e560296
00000804
0736f016
60c3fd96
a2c371c3
105c0070
7c8017a4
32c34c69
0040341c
57546007
75cc58c3
2026002c
36644046
326430c3
4d546007
575c5aac
a81201e9
0404325c
04c4125c
60376c80
8bcc28c3
101c06c3
400600c0
466435c3
465c90c3
7aac17c4
04c4035c
01e9575c
17c7353c
0564165c
2e8c6c80
200751c3
24091654
400620b7
04942027
00415f5c
209725c3
361c31c3
133c0003
313cfff0
12c3f88c
207713a3
00215f5c
0030343c
32835f86
18c36180
0664415c
29c306c3
2ac32980
466435c3
355c58c3
06c30404
366419c3
e0760396
08040f56
60c37016
42c351c3
4006660c
1000211c
67d23283
25d225ac
6ecc622c
366404c3
67d2758c
6dac7a2c
153c04c3
36640300
62f270ec
7fe51004
710c70ef
710f6c0c
712f62f2
6e4c786c
153c06c3
36640040
08040e56
0336f016
60c3ff96
42c391c3
0a352167
301c0116
311c0b84
6c0c0000
366403a6
f10c8056
65f27d8c
9abc04c3
1d8f090e
60061d90
680f28c3
9d8c7a2c
06c3ad8c
273c17c3
343c0040
56640980
323c5d8c
62320980
04d6325c
025c0026
325c04c6
6f9204e4
04e7325c
6d6c7a2c
17c306c3
301c3664
28c30800
865c694f
065c0427
00720a69
2f5c0037
265c0001
393c0a6d
001c100c
011c7300
2c002010
4c000045
808b383c
4026680e
0196440e
0f56c076
00000804
800c1016
200604c3
0004111c
093ceabc
06a4345c
1524335c
345c66f2
60252604
2607345c
08040856
40c31016
0604205c
6492686c
305c686f
6c6c0604
0002341c
02c66bd2
1341145c
087300bc
0604245c
6192686c
0856686f
00000804
40c31016
06a4305c
2580233c
6025688c
68cc688f
28af63f2
2c0f0053
600628cf
0226640f
1341145c
087300bc
145c0226
a2bc1341
08560872
00000804
0136f016
71c360c3
801ca006
383c0001
3783500d
453c6dd2
04c30070
1341165c
087300bc
165c04c3
a2bc1341
a0250872
ee94a187
0f568076
00000804
0136f016
80c3fe96
52c371c3
8146c88c
2954e087
1c94e0a7
21c338eb
000f241c
60777969
00213f5c
42c33064
1b156007
13c36057
007f141c
3f5c2037
796d0001
0010423c
0f358067
fff0423c
01160193
0b84301c
0000311c
001c6c0c
366400ad
80068056
03c7343c
115c18c3
4c8006a4
31c338cb
2000341c
e0876fd2
688c0d54
688f6025
64f268cc
740fa8cf
28ac0073
a8af340f
688c0193
688f6025
63f268cc
0053a8af
a8cfac0f
740f6006
04c380e5
135c38c3
00bc1341
04c30873
135c38c3
a2bc1341
02960872
0f568076
00000804
0136f016
40c3ff96
c5ac51c3
ff60363c
12356027
1054c107
06a4205c
1344325c
325c64f2
68d21524
0070063c
1341145c
08732cbc
e0060a73
0070863c
01c1255c
750c48d2
65f26037
00012f5c
01c5255c
01c1355c
750c63d2
74ac68f2
722c66d2
04c36e6c
366415c3
6007750c
54292054
341c32c3
60070002
722c1a94
04c36e8c
029315c3
07a4345c
100462f2
345c7fe5
345c07a7
6c0c07c4
07c7345c
345c63f2
706c07e7
04c36e4c
36642085
07c4145c
e9942007
6af274ac
68f2750c
0070063c
1341145c
0872b8bc
08c30133
1341145c
0872d0bc
e026e3f2
0196f653
0f568076
00000804
0736f016
40c3ff96
e5ac51c3
273cc50c
60260080
200d833c
0054a01c
2010a11c
007c901c
2010911c
65d274cb
04dc6027
1253000a
0a93245c
374332c3
0001341c
a4dc6007
e0e70009
245c1fb4
40070a61
d50c1b94
01c1355c
265c6df2
323c01e9
245c17c7
6d000564
341c6c0c
60070001
722c2e94
04c36e2c
25c316c3
d50c3664
e994c007
e14704b3
245c2294
40070a61
d50c1e94
40067a0c
0800211c
60073283
265c1654
323c01e9
245c17c7
6d000564
341c6c0c
6bf20001
6e2c722c
16c304c3
366425c3
c007d50c
0053e694
355cc9f2
600701c1
c0065154
01c5655c
700c09b3
045c2c4c
40290544
2894e147
601c7a0c
611c3000
36830008
20946007
04c4345c
60276cc9
323c0894
6580300c
0464335c
14946007
335c706c
204606a4
708c3664
0331245c
3e87023c
40a62c6c
0fe4301c
0000311c
5abc6cac
74290874
60376172
00016f5c
722cd42d
04c36d2c
366415c3
54ce4026
60060233
2ac374ce
39c30811
722c0c11
04c36fac
366415c3
750c05f2
b4dc6007
0196fff5
0f56e076
00000804
3f36f016
50c3f496
105c81c3
22771384
406ca390
38c342b7
cd0c2db0
01c0183c
40062237
01cd235c
305c6006
705c25e7
465c0564
205c01e9
323c0a69
68d20024
41774192
00a14f5c
0a6d405c
1dc33413
32c3440b
640e6025
11a3305c
622c67d2
36646dec
34dc0007
255c0019
323c0a69
6bd20044
41374292
00810f5c
0a6d055c
101c798c
2c0f0201
17c7343c
c384c7c3
0147493c
402681b7
900d323c
316433e3
393c61f7
63120040
133c7580
20f71ac0
03a0493c
355c80b7
602525e4
25e7355c
12dcc007
798c0015
6bf262f7
001c0116
011c0b84
600c0000
00a5001c
80563664
6c1062d7
60077a0c
3b3c3b15
65d20024
01f9265c
34944007
345c8257
001c0a24
011c8000
10c30000
0a5431e4
201c0116
211c0b84
680c0000
36640326
82578056
0a24345c
8000001c
0000011c
31e410c3
201c1794
245c0400
61260a27
09a6355c
06c4355c
0a13145c
3e87013c
40062c0c
0fe4401c
0000411c
5abc70ac
ab3c0874
0ac30024
1f540007
2584255c
01f9165c
13942007
49806197
6025684c
355c684f
60072804
09c32b54
0fe4401c
0000411c
b4bc30cc
04530873
68000197
40254c2c
03934c2f
2804355c
09c369d2
0fe4201c
0000211c
b4bc28cc
355c0873
81972584
680c4e00
680f6025
25a4255c
6025680c
2006680f
20ce0dc3
7a0c206e
211c4006
32830020
15546007
0283365c
900c80d7
00d76e00
2097600f
1e1d253c
34e442c3
01d70814
055c30c3
30830f63
0f66355c
00143b3c
01166af2
0b84101c
0000111c
0346640c
80563664
80043b3c
00046ed2
00040004
00040004
00040004
355c0004
60251964
1967355c
e2d27ac3
762ce026
05c36f0c
27c316c3
365c3664
67320201
400664d2
1495255c
8c6c75ec
17c306c3
35c329c3
7a0c4664
411c8006
34834000
2c546007
0007931c
265c29b4
1cc301f1
07a9415c
324334c3
0001341c
1e546007
0080323c
303c0026
47ec300d
60073283
465c1594
343c01e9
c3c317c7
0564055c
e037c084
6a8562d7
05c36077
26c318c3
fabc3cc3
60c30919
1ac30833
265c25d2
400701f9
762c4094
05c38f8c
26c318c3
46643bc3
345c8297
02170644
366416c3
355c980c
602507a4
07a7355c
07e4355c
655c64f2
005307c7
655ccc0f
000607e7
762c180f
08c36dac
02c01f3c
18c33664
452c650c
48d265d2
66d264ec
44f201d3
68ec28c3
01166ad2
0b84001c
0000011c
0b06600c
80563664
3b3c64c3
60072004
ffeab2dc
000b931c
931c0454
0f940009
70ec48c3
70ac6cf2
05c36af2
111c2006
eabc0004
05c30904
0910dcbc
0c960006
0f56fc76
00000804
0736f016
40c3fa96
62c371c3
a06c93c3
0100af3c
0684355c
40061ac3
29c33664
355c4dd2
04c30684
40261fc3
0f3c3664
1fc30080
f4bc2ac3
611708fc
043436e4
7fe56157
c1376177
69d239c3
1f3c07c3
2f3c0100
0cbc0080
009308fd
4157dc0f
06965c2f
0f56e076
00000804
205c1016
40070a61
305c3454
600711a3
105c3054
27d21253
1283205c
fff0313c
271523e4
1264405c
1f542007
1283205c
602532c3
1286305c
301c0313
311cc350
23c30000
06b442e4
9cbc04c3
80060895
001c0193
011cc350
9cbc0000
301c0895
311c3cb0
9180ffff
e8948007
00b30026
405c8006
00061286
08040856
3f36f016
60c3f996
85b0b1c3
0f63105c
3c4331c3
0014433c
1bc38037
4006a50c
622c44ee
15c36d4c
36642cc3
0243355c
962c6077
160c8177
111c2006
01830800
28540007
01e9155c
17c7313c
265c93c3
92840564
4e9039c3
87d24ac3
1783265c
336431c3
1fb423e4
0a61165c
01162bf2
0b84301c
0000311c
04666c0c
80563664
a65c0253
40060584
01ed255c
0564965c
455c0153
343c0279
a3c30cc7
0584165c
90c3a184
100c3c3c
7300201c
2010211c
41b74d00
7302401c
2010411c
80b78e00
00f70006
0137e026
758cd0c3
0bc36bf2
090eacbc
84dc0007
0bc3001c
090e9abc
7aac158f
2e8c158c
08cb9cbc
2026758c
0636135c
32c3560c
760f6992
455c8057
01570246
2017162f
757224d2
00f3760f
fdff301c
ffdf311c
560f2383
341c760c
5a2c0800
6aac67d2
1cc306c3
36642bc3
15903373
06c3898c
253c15c3
383c0040
46640980
8006760c
4000411c
60073483
c31c5a54
57b40007
01f1255c
415c19c3
34c307a9
341c3243
60070001
07ec4c54
0080323c
14c38026
31c31323
6bf23083
00c7323c
698029c3
07e3235c
0263355c
245423e4
308331e3
63ef09c3
01f1155c
00c7213c
435c6100
323c0813
5aac0fc0
2b8c0180
08cb9cbc
01f1255c
00c7323c
618009c3
0816435c
01f1155c
00c7313c
255c6180
235c0263
455c07e6
343c01f1
321c00c7
06c300fc
49c315c3
345c5180
3ebc07a1
00f7093d
005c08c3
00070633
001332dc
6d6c7a2c
15c306c3
760c3664
0400341c
751c63d2
1bc33000
25d2248b
694c28c3
694f6072
60076117
000fb4dc
80074ac3
0dc32154
1e940007
2006760c
0800111c
6cd23183
71eb578b
0001d01c
12b423e4
60cc0ac3
0024d33c
c31c01b3
08b40009
68cc2ac3
0002341c
0002d01c
d01c63f2
365c0000
6af20a61
88d24dc3
15c306c3
3cc32dc3
090d28bc
355ce372
67320211
e17267d2
28c4365c
365c6025
c31c28c7
1e94000a
17a4165c
4c697480
341c32c3
60070008
760c1554
0100341c
10546007
435c38c3
06c30544
255c362c
b4bc0279
100f090e
345c48c3
00060544
355c0c2f
67320201
46546007
415c18c3
06c30544
255c362c
b4bc0279
100f090e
325c28c3
80060544
055c8c2f
303c0279
a3c30cc7
0584165c
548ca184
345c4ac3
64120653
045c696e
30c30653
33646025
0656345c
0fff331c
40060435
0656245c
760ce772
411c8006
34832000
373c65d2
73c30c05
265c7364
686c0604
0010341c
741c63f2
686cff3f
686f6472
0604265c
6572686c
c31c686f
02940009
101ce672
111c0448
640c2010
0001341c
01166af2
0b84201c
0000211c
0486680c
80563664
6d4c79cc
366406c3
3bc38026
01cd435c
341c762c
6ff20580
09e4365c
0b3561c7
101c0116
111c0b84
640c0000
00a3001c
80563664
684c28c3
000f341c
0400201c
23c362f2
72c327a3
808b383c
700e8097
400e0197
2804065c
20540007
01f9355c
0a04165c
32e421c3
365c1994
2c8c06c4
401c2cc3
411c0fe4
70cc0000
08745abc
011701b3
283c618c
4e4e108c
0253155c
101c21c3
21a38000
455c4e6e
2bc30253
710048eb
236423c3
4cee3bc3
32e46c8b
760c0b14
0200341c
62f240d7
a137540c
52c343d2
0796c673
0f56fc76
00000804
3f36f016
50c3fa96
005c61c3
30c30a93
3043074b
0001341c
155c66d2
20070a61
001a52dc
0448c01c
2010c11c
0b84d01c
0000d11c
e007f8ac
001992dc
28c31c90
275c49e9
38c301ed
06320d29
1f5c0137
175c0081
b55c027d
a55c0584
475c0564
935c01e9
79ac0021
e4dc6147
746c0010
142c6dcc
40462026
30c33664
69f23264
033c79ac
155c0070
2cbc1341
2dd30873
6007790c
0016b4dc
62f2788c
7fe51004
78ac788f
78af6c0c
78cf62f2
333c79ac
055c0147
4c002584
6025686c
255c686f
684c25a4
684f6025
2384255c
18c37500
135c2449
323c23a5
40062420
371d253c
6c4938c3
10546007
17c305c3
09019abc
e0f7f8ac
c4dce007
740c000b
00610f5c
0ab5035c
1cc316b3
341c640c
60070001
7e0c1054
211c4006
32830800
19546007
17c7343c
61810ac3
0001341c
11946007
341c7e0c
66d20040
155c0066
00bc1341
746c0873
05c36e4c
0040173c
12133664
5c8c19c3
56ac6500
04c4025c
64092c00
00d0331c
01172f94
0cc7303c
69a22bc3
10946027
0644355c
341c6c0c
6ad20010
233c31c3
02c3009e
00b70472
00412f5c
67094c0d
16946067
40074729
075c1394
303c01e9
055c17c7
4c000564
30c30769
003c341c
65856232
359d323c
315c6412
762c00fe
05c38cac
26c317c3
466439c3
2384355c
2420233c
2c0b7c8c
271d153c
686828c3
39156007
0149165c
011627f2
680c2dc3
36640306
796c8056
0149065c
3fe510c3
2f5c2077
41770021
00a10f5c
014d065c
2a1d133c
5e0c3daf
7b7232c3
08c37e0f
31c320cb
1000341c
60066dd2
4800311c
5e0f23a3
243221c9
2f5c2037
275c0001
762c01f5
05c36eec
5dac17c3
7e0c3664
7e0f7c72
602578ec
792c78ef
f90f63f2
ec0f0053
6006f92f
355c7c0f
60252384
2387355c
d9dc61e7
0006ffed
2387055c
18c3db13
32c34449
0001341c
365c65d2
60070149
788c6954
100462f2
788f7fe5
6c0c78ac
62f278af
79ac78cf
0147333c
2584055c
686c4c00
686f6025
60e779ac
275c1cb4
323c01e9
055c17c7
6c000564
341c6c0c
60070001
155c1094
2df20a61
6e4c746c
173c05c3
36640040
1944355c
355c6025
d3b31947
8cac762c
17c305c3
39c326c3
762c4664
05c38fcc
26c317c3
466438c3
11a3355c
b4dc6027
255cffe8
40271233
ffe864dc
1243755c
7fe537c3
12a4455c
055c39ac
43e40a93
323c0b94
33e3100d
355c3083
00060a96
12a7055c
323c0173
30a3100d
0a96355c
0010343c
12a7355c
0696ccd3
0f56fc76
00000804
105c1016
313c1471
405c17c7
2e000564
315c6006
315c0ae7
315c0b07
315c0b27
23640b47
0b76215c
03f0323c
0b86315c
fc00323c
0fff341c
0b66315c
08040856
400b1016
802b6520
341c6e00
4026001f
300d323c
204c33e3
604f3183
800b0193
602534c3
0fff341c
313c600e
341c0010
602e001f
604b202b
075431e4
100d323c
3483804c
ec546007
08040856
400b3016
133c6520
402bfff4
433c6500
602601f4
a04c3423
604f35a3
7520a04b
001f341c
061413e4
0010343c
001f341c
0c56604e
00000804
402c1016
0e9421e4
62f2600c
7fe51004
602c600f
602f6c0c
12946007
0213604f
680c23c3
045431e4
23c37cf2
640c0073
680c680f
404f62f2
7fe5600c
0856600f
00000804
0136f016
41c350c3
83c372c3
68d2658c
6dac622c
260502c3
40063664
720c518f
211c4006
32831000
762c66d2
07c36ecc
366431ac
0263645c
16c308c3
09191ebc
335c746c
073c0644
14c301c0
355c3664
602507a4
07a7355c
07e4355c
455c64f2
005307c7
455c8c0f
600607e7
28c3700f
36e4680b
363c0794
341c0010
28c30fff
8076680e
08040f56
100c213c
322361e6
205c33e3
328307c4
07c7305c
00000804
22121016
312361e6
405c33e3
348307c4
21234372
305c32a3
085607c7
00000804
40c33016
4fd251c3
100c313c
07c4205c
308d323c
0074233c
5fe546d2
d2bc44d2
00b30919
15c304c3
0919c6bc
08040c56
3f36f016
60c3fc96
52c32037
01e4af5c
025c2417
203c01f1
221c00c7
4d0000fc
558c4077
0633925c
60b7682c
0000801c
c01cd8c3
4ac30001
052b8ef2
208c803c
0140d13c
02e3465c
840934c3
33c43403
f88cc33c
0980123c
e00620f7
355c7410
4ac30263
40072cc3
4ac31994
14948007
233c38a4
1accfff4
21e410c3
1ac30d34
341c4552
8026001f
300d343c
403c0dc3
34832a1d
202662f2
e7d241c3
6dcc7a2c
15c306c3
366424c3
155c85d2
200701f9
760c1494
211c4006
32830100
7a2c67d2
06c36e0c
409715c3
06c33664
401715c3
82bc6057
01730919
0540153c
20d7e2f2
6006446c
680b640e
680e6b72
fff0393c
936493c3
04d209c3
5bc3e025
0bc3f613
fc760496
08040f56
40c33016
036403c3
18542007
22f22232
323c2026
201c00f4
211cc950
523c0011
313c399d
133c528d
01e4188c
64200734
0303545c
0350141d
00060053
08040c56
0136f016
313c62c3
205c17c7
ad000564
0b63855c
59a038c3
fff4323c
05dc6fe7
65320009
0570733c
7a1d453c
01f4323c
323c4026
13c3300d
02c31483
d4dc2007
34a30008
7b9d353c
0b73355c
63e401c3
000844dc
0b24355c
1b947fe7
0b04255c
0ae7255c
0b07355c
0b44355c
0b27355c
0b47155c
0200363c
0b76355c
0b83755c
640537c3
0b86355c
0200383c
0b66355c
0b24355c
0b04155c
1d947fe7
0ae7155c
0b07355c
0b44355c
0b27355c
755ce006
155c0b47
31c30b73
355c6405
255c0b76
32c30b83
355c6405
755c0b86
37c30b63
06736405
333c33e3
433c080d
053c0b8d
255c15c0
34c30ae4
089326bc
34236026
155c7fe5
31830b24
4a204406
255c3223
32a30b04
0b07355c
1640053c
0b44155c
0b24255c
26bc34c3
24c30893
755c2364
6b800b73
0b76355c
0b83155c
355c6880
755c0b86
6b800b63
0b66355c
263c01b3
622c0010
241c6c2c
36640fff
0b04355c
355c7f72
00060b07
0f568076
00000804
42c3f016
0564605c
01e9215c
0279515c
0cc7353c
0584705c
660caf80
0002341c
17546007
05c4255c
0804323c
7f546007
2a0b023c
02e0153c
a00632c3
4000511c
523c3583
6007144b
523c1954
02d3138b
17c7323c
323c5981
60070024
023c6854
153c288b
32c302e0
711ce006
37838000
164b523c
523c63d2
0147158b
02073354
00271854
640c4d94
640f6025
31c367f2
023e033c
402520c3
440b4c0e
353c500e
6d72700c
642b702e
a44b704e
07f3b06e
6025640c
67f2640f
733c31c3
27c3023e
4c0e4025
0006b00e
440b102e
642b504e
a44b706e
10aeb08e
10ee10ce
112e110e
640c04d3
640f6025
31c367f2
023e733c
402527c3
640b4c0e
408c233c
5f00341c
32c323a3
700e6d72
700c353c
04096d72
702e30a3
504e442b
706e644b
640b0113
6025700e
353c640e
702e700c
08040f56
3f36f016
a0c3f296
52c341c3
0279015c
0cc7303c
115c1ac3
0c800584
32c3520c
711ce006
37830800
69d263c3
01e9145c
17c7313c
775c7ac3
cf800564
6e7232c3
145c720f
223701f1
225c2ac3
47f20a61
335c3ac3
345c0a01
009301fd
745ce026
508c01fd
1f3c6006
ed6202c0
6045e5c1
fc946187
60276009
60670354
b63c0d94
c01c0480
20060100
3f3c2277
62b70320
02c0df3c
203c0193
42b70080
0000c01c
0200701c
b1c3e277
0320df3c
440b1bc3
341c32c3
520c0001
18546007
617232c3
305c720f
233c05c4
133c0804
601c2a0b
43f24000
12c362c3
345c6006
e00601ed
0266745c
0000901c
32c30493
111c2006
31834000
f4dc6007
103c000e
205c0b40
93c305a3
0266245c
32c3440b
341c6025
640e0fff
323c580c
69d20024
341c720c
123c0010
601c288b
63f24000
16c3c006
e006720c
0004711c
801c3783
62f22000
034683c3
701c01f7
29c30080
630644f2
79c361f7
30c301d7
03c37f45
c0070364
21471354
42460754
05542207
20274086
41060294
250021d7
3f5c21b7
61f700c1
03c36100
20060364
306e304e
201c704c
211c00ff
32839fff
704f7f92
00e13f5c
704c710d
6c0b233c
323c4100
704f6c1b
305c0ac3
6c0c0644
0010341c
1000201c
23c362f2
c1a32257
63723cc3
03a306c3
78a380a3
540e27a3
342e2006
480b2bc3
3bc3544e
746e6c2b
fc4b7bc3
0297f48e
14ae000b
242b2297
429734ce
54ee484b
6c0b3dc3
7dc3750e
f52efc2b
004b0dc3
345c154e
64120263
6186756e
200719c3
320c1654
400631c3
0200211c
42063283
23c362f2
311c6006
13830040
22f26406
e21731c3
32a327a3
61a6758e
6112c7d2
14c30ac3
4ebc5580
01d7091b
606530c3
233c6132
1ac30fe4
27c1315c
0010023c
60270037
301c1994
353caaaa
3f5c271d
e0660001
371d753c
0010133c
3f5c2177
201c00a1
253c9640
033c371d
01370010
00813f5c
101c0473
153caaaa
3f5c271d
40660001
371d253c
0010033c
3f5c00f7
20060061
371d153c
0010733c
3f5ce0b7
01930041
23c36217
323c4585
3980080c
259d263c
0001901c
3264e1d3
0ac32006
27c5105c
080c733c
0f5ce077
045c0021
218601dd
01e5145c
fc760e96
08040f56
0006600c
1341135c
0872a2bc
00000804
0f36f016
90c3ff96
6010c32c
0ba4a05c
0704305c
0003835c
0ac3ec2b
b3a0802c
2bc305c3
17a4125c
08cb9cbc
213c300c
323c230b
67d20084
0007241c
323c31c3
700f231b
64327029
0f5c6037
055c0001
19c301d5
700c46ec
0fff341c
6e008b0c
0006778e
178b160f
67a018c3
023530e4
73c330c3
f4ce7364
6c2c3ac3
c047748f
40060694
44af1ac3
02b346c3
c0c78026
1a3c1294
642c0100
1ff0233c
702c4ac3
01ff321c
301c2303
2383fe00
43f28006
8046442f
1ac34006
63a0442f
836483c3
200c343c
733c6580
c0260040
08c30493
336438c3
0200331c
001c0335
03640200
088c263c
0014163c
0067323c
60c56c80
371d053c
0037323c
60856c80
253c5c0c
60063b9d
087f373c
642018c3
836483c3
c0258025
600738c3
343cdb94
4ac3200c
433c7180
03b30040
088c263c
0014163c
0067323c
60c56c80
053c0006
323c371d
6c800037
20066085
3b9d153c
27d2300c
40060bc3
08e6e6bc
500f4006
8205c025
e335c0a7
445c49c3
87d20361
62cc09c3
15c36ccc
08333664
01d1155c
19942007
325c29c3
602507a4
07a7325c
07e4325c
525c64f2
005307c7
39c3ac0f
07e7535c
940f8006
00a66c4c
a2bc2c0c
04b30872
78bc0e06
201c08cc
211c0b1c
680c0000
680f6025
63f2684c
0053a82f
301cac0f
311c0b1c
ac4f0000
140f0006
82bc0e06
004608cc
125c2bc3
301c1341
311c0fe4
4d0c0000
08c8d4bc
f0760196
08040f56
0136f016
a32c72c3
0293615c
0f94a047
32c3440b
1f866065
640e3083
27c301c3
363c8006
833c0010
0213180c
f794a027
30c3040b
00ff321c
ff00201c
fdd33283
680f600c
684e604b
81054105
48e40105
a047f894
363c1094
5d80180c
080c363c
013c6025
30c3399d
3f866065
325c3183
0293ffe6
1294a027
080c363c
313c6025
201c399d
331c0200
03b40100
0100201c
180c363c
235c7d80
363cffe6
1d80180c
0f568076
00000804
0336f016
e00c40c3
93c36e24
305cf524
835c0764
a0060021
0edc601c
0000611c
382c02f3
62f2780c
7fe51004
642c780f
62f2782f
345c784f
64d20361
6acc502c
7c6c7ff2
05a4335c
366407c3
58e4a025
393ce994
62d24004
c076f324
08040f56
3f36f016
60c3fc96
92c3d1c3
4010c3c3
20b7232c
0764205c
305c4077
001c03f9
011c0edc
60070000
8e241d54
1ac3f524
135c66ac
9cbc04e4
409708cb
608732c3
78ac0794
301c4c2c
0c0c0b00
20062664
03fd165c
4004343c
42dc6007
f3240008
a02c1033
7e54a007
680f29c3
60f783c3
73c360d7
365ce025
73e403f1
340b45b4
01162af2
0b84201c
0000211c
0246680c
80563664
0000b01c
0283355c
80d767f2
202714c3
b01c31b4
40970001
602732c3
940b1494
321c34c3
685200ff
365c8384
83e40da3
01160a35
0b84201c
0000211c
0226680c
80563664
6c2c79ec
06c36037
2dc315c3
00614f5c
801734c3
d0c34664
640c19c3
6d00540b
b42c640f
3bc3a6d2
e0f764f2
e0d7f6d3
f02f8057
0894e027
325c2ac3
4c4c18a4
4c4f4025
365c01f3
4ac303f1
18a4245c
059473e4
6025680c
0093680f
6025682c
301c682f
311c0edc
6c2c0000
0283235c
323c4ad2
6027ffc0
406606b4
440f1cc3
00b30026
4c0f3cc3
0006ff93
fc760496
08040f56
fe96f016
51c340c3
40072364
606c1854
40271fc3
335c0e94
40060684
1f3c3664
00060040
711ce006
6f3c8000
03b3ffc0
0524335c
14c30fc3
fe533664
0b64305c
605c6037
c0770b84
0112fd73
208d373c
62d23483
50e40072
02a002b4
44074025
3f85f594
045416e4
4006840c
0296fdf3
08040f56
800cf016
345cf1cc
633c06a4
b90c1e00
1c54a007
6dac70cc
366404c3
7322301c
2010311c
4c0e4006
7320301c
2010311c
6c0c4c0e
70cc66d2
04c36d8c
00d33664
04c37c6c
25c316c3
0f563664
00000804
200c3016
0544315c
66126c29
0580533c
215c804c
680c0624
680f6025
6c4c65cc
328001c3
0c563664
00000804
0f36f016
40c3ff96
705c81c3
a05c1824
505c0664
305c1544
53e40353
145c1635
29d21481
1864345c
345c6025
40061867
1485245c
1864345c
0a356067
0343545c
045c0086
00931867
145c2006
345c1867
2ea00b64
0b84245c
023435e4
345c5fe5
67f212e4
9000001c
0001011c
12e7045c
1323345c
c02666f2
1326645c
1336345c
1333645c
12e4045c
0037303c
53e46232
24000535
023410e4
38c34025
24002c30
10e4a006
40250234
fff0363c
645cc5f2
36c31323
63c37fe5
92e46364
92e40714
38c31494
b1e46c10
08c31034
6420000c
1887345c
12e4145c
32e421c3
301c0f35
345c03e8
01531887
a8072400
353c0654
53c30010
fad35364
0026c026
3da90037
1d8927d2
0b0d303c
7f327fe5
1f5c6037
3ac30001
32c34c0c
ffe0001c
0001011c
60073083
40261794
1ac323d2
545c458b
345c1884
60271521
323c18b4
045cfff0
333c1323
6f00028d
12e4145c
128d333c
545c0173
29d21884
614b323c
245c7fe5
333c12e4
b580228d
7d8d6026
68c37dad
7700d80c
706c7c0f
0524335c
14c308c3
18c33664
345c040c
6c0c1824
033530e4
ac207c0c
05c3bc4f
f0760196
08040f56
40c31016
23c302c3
341c70ec
68d20001
7172640c
600c640f
600f6072
680c0093
680f7072
341c70ec
68d20002
7572640c
600c640f
600f6172
680c0093
680f7472
341c70ec
68d20004
7d72640c
600c640f
600f6372
680c0093
680f7c72
341c70ec
68d20008
7972640c
600c640f
600f6272
680c0093
680f7872
08040856
40c31016
eabc3fe6
0286093c
1341145c
087300bc
08040856
698cff96
0201201c
64294c0f
241c23c3
403700fd
00013f5c
65ac642d
1341205c
0070033c
00bc12c3
01960873
00000804
0f36f016
40c3fe96
605c91c3
705c0604
60700544
04c4805c
02c64010
1341145c
0872d0bc
323c586c
66f20014
13a1345c
e4dc6027
345c0012
ac091504
4d54a007
0104323c
66f2a006
6c4c710c
366404c3
586c50c3
0104323c
15946007
644918c3
05946027
31c3382c
0d3553e4
13a1345c
33946027
1384345c
0a13135c
3e87313c
2bb453e4
65ac19c3
27b46027
0044523c
1f94a007
08bc301c
2010311c
1bc3ac0f
04c365ac
0ef0101c
28c33664
60276849
545c0494
00f30aa6
13a1345c
06946027
0ab6545c
c4bc04c3
786c0901
786f6272
6172786c
1c33786f
323c586c
60070044
28c36b54
60276849
145c0994
31c30aa3
0eff351c
0aa6345c
345c0193
602713a1
045c0b94
30c30ab3
0aff351c
0ab6345c
c4bc04c3
786c0901
786f6372
644918c3
0d946027
61ac09c3
04b46027
5580784c
09c30253
101c41cc
03730400
13a1345c
0b946027
1384345c
0a13235c
3e87323c
4c00184c
01b32006
301c0116
311c0b84
6c0c0000
00d3001c
80563664
12c34006
618c0bc3
366404c3
65ac19c3
16356027
ac4938c3
1294a027
001c71cc
2c8c012c
301c4206
311c0fe4
6cac0000
0874c4bc
722c301c
2010311c
345cac0e
4c4c0624
4c4f4025
323c0e53
60070084
345c6e94
2c091504
51542007
284928c3
09942027
61ac09c3
49b46027
03c3782c
453550e4
13a1245c
09944027
1384345c
0a13035c
3e87303c
393553e4
1e942027
f060001c
7c6f7400
08958ebc
60803c6c
7c697c8f
61723264
2f5c6037
5c6d0001
32647c69
60776572
00213f5c
0ac37c6d
6c2c60ec
366417c3
40270353
716c1894
05c36cec
366414c3
11940007
684928c3
04946027
0aa6045c
345c00f3
602713a1
045c0694
04c30ab6
0901c4bc
604908c3
05946027
6d0c71ec
366404c3
08bc301c
2010311c
4c0f4006
145c0066
00bc1341
02c60873
1341145c
0872b8bc
f0760296
08040f56
40c31016
145c02c6
48bc1341
00070873
245c1094
686c0604
686f6272
145c02c6
a2bc1341
02c60872
1341145c
087300bc
08040856
40c31016
0664105c
6ef2648c
6cf264ac
001c640c
011cffe0
30830001
458b65f2
602643f2
048c658e
44ac05f2
36944007
440c07d3
616b223c
345c440f
600712e4
0a121054
01a00133
233c640c
4025614b
615b323c
345c640f
03e412e4
04f3f534
402632c3
615b323c
0433640f
12e4345c
11546007
00d34a12
058b49a0
602530c3
345c658e
045c1323
333c12e4
23e4028d
01b3f434
458e4026
640c0153
615b303c
058e640f
1323345c
fc3376d2
08040856
0136f016
60c3ff96
0664405c
705c0210
648c0644
540ba980
323c700c
700f081b
4832540b
105b323c
542b700f
10db323c
233c700f
40370014
73544007
0018341c
1469205c
0e946107
01164ad2
0b84301c
0000311c
01466c0c
80563664
536d4026
4af201b3
301c0116
311c0b84
6c0c0000
36640166
60468056
700c736d
323c544b
700f615b
304e346b
706f748b
323c54ab
333c81ac
706f3e87
111c2006
21c37fff
023532e4
350b306f
352b21c3
812c313c
554b708f
556b12c3
80ac323c
758b70af
35c3718e
063e133c
213c502c
502f0c1b
68326c0b
00f4133c
313c32c3
702f24db
213c5c0c
5c0f201b
00f4323c
32c369d2
323c41e6
7c0f201b
7092702c
35c9702f
3e87313c
28c3704f
06c3680c
18c33664
06c3644c
366414c3
6c2c79ac
00f306c3
00012f5c
1525205c
648c18c3
00263664
80760196
08040f56
0336f016
70c3ff96
c00c81c3
0644565c
0544405c
233c640c
4037104b
00013f5c
165c704d
20070361
74091494
05946027
13c36017
20542027
40067429
1d946027
32c34017
0002361c
233c7fe5
02b3f88c
4e6c782c
6127680c
60670354
41060394
61470193
60870354
201c0494
00b30200
402668ec
444662f2
0c6c38c3
945c106f
2c0c0011
0001931c
313c2194
61070184
07f20694
607232c3
0213714e
04946207
637232c3
0116ff53
0b84301c
0000311c
001c6c0c
366400b7
7b2c8056
60277f85
714b16b4
714e6072
313c0253
61070184
0af20994
31c33429
0001341c
518e65d2
620700d3
32c30494
718e6372
6c6c7e0c
18c307c3
78ec3664
184c6d0c
366414c3
c0760196
08040f56
40c37016
0664605c
205ca20c
680c0644
202b333c
74ac680f
744c3664
16c304c3
71ac3664
04c36c2c
0e563664
00000804
005c42ac
290c0664
08cb9cbc
00000804
40cb6006
602548f2
03946187
00930026
ff130785
08040006
323c440c
60070104
323c1354
68d200f4
1004323c
32c365d2
640f6572
440c046f
00f4323c
32c365f2
640f6572
0804046f
40c31016
280c01c3
0104313c
313c69d2
62f200f4
680c05d2
680f6672
0856884f
00000804
0336f016
63c390c3
726471c3
836482c3
58cb583c
423c4049
6dec0fe4
06c36ccc
0014123c
54e43664
343c1714
6f80ffc0
12b453e4
2006f9ec
49c37620
383c5180
00260074
300d303c
34838869
10c362d2
06c37cac
c0763664
08040f56
400c10c3
6c2c68ec
115c02c3
36640544
00000804
50c33016
734c806c
60263664
730c07f2
366405c3
002602d2
03c330c3
08040c56
604c4006
6ca0206c
021532e4
02c34026
00000804
0644205c
680c25d2
67927072
0804680f
c1ac7016
0644505c
2007540c
32c31054
740f7272
2724005c
408638ec
0fe4301c
0000311c
c4bc6cac
02130874
200632c3
0004111c
6ad23183
1333105c
32c327f2
0c9b313c
78cc740f
0e563664
00000804
405c1016
0f260544
08cc78bc
2a4c534c
10096026
33e33023
6a4f3183
82bc0f26
085608cc
00000804
40c31016
6fac606c
00073664
445c1094
0f260544
08cc78bc
464c334c
10096026
32a33023
0f26664f
08cc82bc
08040856
002630c3
0989235c
002648d2
1341135c
087348bc
002602d2
00000804
005c30c3
135c16a4
56bc1341
02d20873
08040026
40c31016
0a93205c
3a8c323c
245c03c3
02831684
1341145c
087356bc
18940007
1384345c
09c3235c
341c32c3
65f20002
335c700c
6cf20584
6eac706c
06a4045c
303c3664
7fe50b0d
f88c033c
00260053
08040856
0136f016
63c350c3
435c0db0
620c0644
011c0006
30830800
72dc6007
40670009
41470435
000924dc
736471c3
155ce5d2
200701f9
500c6694
000632c3
0400011c
6dd23083
7a9232c3
18c3700f
06c364cc
02863664
1341165c
087300bc
341c700c
61e7000f
68f20654
341c760c
64d22000
6992700c
500c700f
341c32c3
60074000
e5d24054
01f9355c
3b946007
341c760c
60070040
32c33654
2000341c
31546007
6a92700c
4e9223c3
323c500f
60070104
00062354
32c3104e
79926c72
780c700f
0744335c
0261135c
135c01c3
213c0269
035c402c
203c0271
135c812c
013c0279
28c3c12c
408628ec
0fe4301c
0000311c
c4bc6cac
02860874
1341165c
087300bc
341c760c
62d22000
700ce4f2
700f7492
323c500c
60070104
323c1854
61e700f4
60070754
760c1294
2000341c
79ec6ed2
360c558c
082c6c4c
0b4b113c
366424c3
6c0c79ec
366406c3
0f568076
00000804
0136f016
e1ac60c3
405c01f0
500c0644
0604323c
1c946807
717232c3
005c700f
3cec2704
301c4086
311c0fe4
6cac0000
0874c4bc
165c0286
00bc1341
500c0873
00f4323c
049461e7
709232c3
700c700f
0060341c
5c946c07
165c0286
00bc1341
500c0873
200632c3
0080111c
63d23183
083332c3
00f4523c
0654a1e7
08f4323c
0080331c
28c32494
04c3698c
50c33664
07d2700c
700f7192
06c37ccc
07133664
700f7172
2704065c
40863cec
0fe4301c
0000311c
c4bc6cac
500c0874
00f4323c
269461e7
353c32c3
02730c1b
2094a007
698c28c3
366404c3
0dd2700c
253c23c3
500f0c1b
2004323c
12946007
707232c3
01d3700f
700f7172
2704065c
40863cec
0fe4301c
0000311c
c4bc6cac
80760874
08040f56
0f36f016
50c3fe96
61d041c3
e00c4070
805c21b0
605c0664
780c0644
323c4026
780f155b
155c0286
a2bc1341
02860872
1341155c
087300bc
0544355c
123c4c69
20770f54
00212f5c
60064c6d
098d355c
0fa4355c
10546007
06c4355c
1604055c
40062c2c
8000211c
0fe4301c
0000311c
5abc6cec
075c0874
05f20361
678c1ac3
366405c3
17548007
6b72780c
355c780f
001c1521
60272710
001c0335
39c33a98
40862cec
0fe4301c
0000311c
c4bc6cac
12530874
0624375c
10c30e49
00f8141c
2f5c2037
4e4d0001
6d6c74cc
366407c3
0361375c
18546007
1114401c
0000411c
680c500c
035c6c0c
0a123653
41262bcc
0fe4301c
0000311c
5abc6cac
700c0874
05c4335c
6d063664
2010311c
0c0f1fe6
0ce4255c
4c0f6285
1ac30c0f
0504315c
366405c3
0361175c
12542007
680c28c3
0018341c
0c946107
6c4c7c4c
0003341c
46546007
6c8c760c
366405c3
28c30833
341c680c
62070018
580c3b94
8004323c
355c6ad2
001c1521
60272710
001c2735
04933a98
602c08c3
011c0006
30830001
323c67f2
6ad200f4
684c28c3
09c367d2
0026604c
366415c3
20070373
301c1954
311c015d
6c0c4130
0002341c
10546007
7a72780c
055c780f
29c32704
408628ec
0fe4301c
0000311c
c4bc6cac
0bc30874
05c360ac
02963664
0f56f076
00000804
40c37016
0664205c
0644505c
0989305c
600703c3
680c2854
0018341c
20946207
08958ebc
245c60c3
323c1471
245c17c7
6d000564
341c6c0c
6bd20001
0c73245c
341c32c3
65d20010
08958ebc
15a7045c
7920548c
04746007
6b72740c
740c740f
0acb033c
08040e56
3f36f016
50c3fa96
09c32010
0644a05c
04c4b55c
9570b470
20cc15d0
655c2177
755c0644
255c0664
44121341
0fe4301c
0000311c
6a008c0c
780c6c0c
66926592
001c780f
011c0b30
23060000
08c986bc
0544355c
123c4c69
20370fd4
00012f5c
7c0c4c6d
0018341c
44946107
0544355c
0c6f1c6c
288c2ac3
0544255c
13e4686c
6ca00334
355c686f
6c6c0544
11546007
08958ebc
0544255c
6080286c
255c688f
68690544
61723264
3f5c6077
686d0021
155c0286
b8bc1341
355c0872
6dac0544
538c8157
133c140c
2664424b
6dcc75ec
366405c3
4046780c
155b323c
0026780f
098d055c
115c19c3
20070361
0013d4dc
255c2713
40071469
001372dc
0544455c
60ec08c3
366405c3
355c106f
0c6c0544
648c1ac3
071430e4
6d6c75ec
202605c3
24533664
70494bc3
4e946027
42bc05c3
75ec08fd
05c36d0c
355c3664
60270981
001134dc
0544455c
60ec08c3
366405c3
155c106f
446c0544
708c4ac3
1b58321c
2d3523e4
1521355c
05356027
ec78001c
646f6800
0544255c
1ac3686c
6ca0248c
8ebc686f
255c0895
886c0544
688f6200
0544255c
32646869
60b76172
00410f5c
255c086d
68690544
65723264
1f5c60f7
286d0061
6dcc75ec
366405c3
04c4355c
4c2d4026
4cc31a33
15c370ec
00073664
000cb4dc
341c7c0c
60070001
000c52dc
632c0dc3
366405c3
0544455c
64ec18c3
366405c3
355c106f
60271521
255c0a35
686c0544
1388331c
321c0435
686fec78
08958ebc
155c188f
313c1471
255c17c7
6d000564
341c6c0c
6fd20001
0c73455c
341c34c3
69d20010
15c4155c
255c6080
6d2015a4
15c7355c
0544355c
988c6c6c
388f2e00
305c09c3
435c0744
04c30281
0289435c
402c243c
0291035c
812c203c
0299435c
c12c343c
0ac365a0
6c20008c
5c4c788f
12544007
341c780c
67f2000f
20067c2c
0001111c
68d23183
0544355c
04c38c6c
023420e4
2ac34c6f
255c288c
686c0544
033413e4
686f6ca0
005c09c3
00070361
01261154
0fe4301c
0000311c
b4bc2cac
301c0873
311c1114
6c0c0000
05e4335c
8ebc3664
255c0895
286c0544
688f6080
0544255c
32646869
61376172
00813f5c
0286686d
1341155c
0872b8bc
445c49c3
8af20ca1
0544355c
01576dac
140c438c
424b133c
75ec2664
05c36dcc
780c3664
323c4046
780f155b
155c2026
355c098d
69d20fa4
301c0006
311c0fe4
2cec0000
0873b4bc
225c29c3
44f20361
28bc05c3
06960925
0f56fc76
00000804
0336f016
845c800c
700c0644
b06cec4c
04c4945c
0286d1ec
1341145c
0872d0bc
0664345c
341c6c0c
61070018
770c0b94
366404c3
40940007
04c3772c
774c3664
07c30693
0544145c
08802cbc
34540027
04c3788c
18c33664
341c640c
60070010
78ec3054
366404c3
4c0c38c3
101c32c3
111c1e00
31830017
23946007
0981345c
1f546007
0644345c
20066c0c
0400111c
60073183
19c31694
60276449
32c30954
4000341c
776c69f2
366404c3
794c05f2
366404c3
028600d3
1341145c
08732cbc
0f56c076
00000804
40c37016
0644505c
32c3540c
111c2006
31830001
35546007
600612c3
0008311c
32c31383
20077092
606c2b94
002c6dcc
36644046
326430c3
028667f2
1341145c
08732cbc
740c03d3
00f4633c
c8f2706c
0564335c
2000001c
366414c3
6f0c01b3
366404c3
0df260c3
206604c3
211c4006
debc0001
740c092e
363c6972
740f0c1b
08040e56
40c33016
0644505c
32c3540c
4400341c
4000331c
32c32294
2000341c
606c67f2
36646eec
6d72740c
706c740f
102c6dcc
40462006
30c33664
67f23264
145c0286
2cbc1341
01330873
206604c3
debc4806
740c092e
740f6a72
08040c56
81ac3016
0664305c
341c6c0c
205c0001
a80904c4
205c35a3
125c1384
31a30bd1
706c63d2
708c0053
0c563664
00000804
fe96f016
a00c70c3
0644655c
001c780c
011cffff
3083fff9
780f7a92
0800341c
47546007
04c4355c
31c32ce9
0001341c
17546007
08958ebc
06e4355c
42208c8c
1583355c
12e4055c
028d333c
091423e4
4006746c
8dec4037
218605c3
466432c3
1521355c
802543c3
0f5c8077
055c0021
175c1525
20070361
101c1954
111c1114
640c0000
6c0c6c0c
4523435c
402524c3
235c2364
035c4526
40c349c4
067424e4
6fcc640c
200607c3
780c3664
780f6b92
6c92780c
0286780f
1341155c
087300bc
0f560296
00000804
41c31016
0644115c
323c440c
6cd20104
707232c3
32c303f2
640f7372
145c0286
00bc1341
08560873
00000804
0644305c
201c6c0c
211c1000
32830406
008669f2
0fe4301c
0000311c
b4bc2cac
08040873
41c37016
0644115c
545cd1ac
440c2724
0104323c
18546007
32c309f2
0c9b303c
78cc640f
366404c3
32c301f3
640f7272
036405c3
408638ec
0fe4301c
0000311c
c4bc6cac
02860874
1341145c
087300bc
08040e56
40c33016
0644505c
6c0c61ac
245c3664
323c1471
245c17c7
6d000564
341c6c0c
60070001
345c1c54
60071469
740c1854
740f6e72
2000341c
706c68f2
04c36eec
740c3664
740f6d72
145c0286
a2bc1341
02860872
1341145c
087300bc
08040c56
40c33016
0644505c
0664305c
341c6c0c
61070018
02860b94
1341145c
0872a2bc
145c0286
00bc1341
245c0873
40071469
740c2454
0104233c
15944007
4010351c
7bff101c
ffff111c
323c3183
740f0b5b
2000341c
706c68f2
04c36eec
740c3664
740f6d72
145c0286
a2bc1341
02860872
1341145c
087300bc
08040c56
40c31016
005c62ac
2d2c0644
08cb9cbc
6ccc71ac
366404c3
145c0286
b8bc1341
02860872
1341145c
087300bc
3fe604c3
093ceabc
6d4c71cc
366404c3
6cac71cc
366404c3
08040856
40c3f016
c26ce00c
205ca06c
45d22753
2784305c
36646c0c
04c3782c
355c3664
04c304a4
355c3664
04c304c4
784c3664
366404c3
ff81301c
0087311c
0361275c
301c45f2
311cff81
345c0007
62861687
16a7345c
0e240116
000b051c
80560f24
111c21e6
275c0182
44f20361
111c21e6
04c30102
0904e4bc
0361375c
786c64f2
366404c3
08040f56
4e2c600c
03c34a4c
06a4135c
08042664
4e2c600c
06a4135c
03c34a4c
26642785
00000804
4e2c600c
06a4135c
03c34a4c
26642f05
00000804
4e2c600c
06a4135c
03c34a4c
00b4121c
08042664
4e2c600c
06a4135c
03c34a4c
00f0121c
08042664
4e2c600c
06a4135c
03c34a4c
012c121c
08042664
4e2c600c
06a4135c
03c34a4c
0168121c
08042664
4e2c600c
06a4135c
03c34a4c
01a4121c
08042664
4e2c600c
06a4135c
03c34a4c
01e0121c
08042664
4e2c600c
06a4135c
03c34a4c
021c121c
08042664
4e2c600c
06a4135c
03c34a4c
0258121c
08042664
4e2c600c
06a4135c
03c34a4c
0294121c
08042664
6c6c62cc
08043664
03c3600c
0b08101c
0000111c
1000233c
093968bc
00000804
101c000c
111c0b1c
ccbc0000
0804092c
fe963016
a00c40c3
72f0301c
2010311c
305c6c0b
75cc0926
05c36d0c
75cc3664
05e4245c
20372026
20772206
05c38d4c
7400101c
2010111c
009a221c
0100301c
02964664
08040c56
2300101c
311c6086
2c0f2010
60854006
60854c0f
60854c0f
60852c0f
60854c0f
08044c0f
60c37016
0e0641c3
08cc78bc
a007b02c
700c1654
100462f2
700f7fe5
6c0c702c
62f2702f
0e06704f
08cc82bc
6c0c7a2c
155c06c3
25c301d1
fcd33664
165c05c3
b8bc1341
0e060872
08cc82bc
08040e56
60c37016
06a4505c
150c8006
620c0313
211c4006
32831000
41ac63d2
408c0053
0644365c
341c6c0c
280b0010
31c364d2
00736c72
6c9231c3
000c680e
e8940007
80878025
a7850354
0e56fc33
00000804
2524205c
105c282c
40061447
148d205c
00000804
800c3016
0624205c
0544345c
101c6dac
111cfe00
31830001
105431e4
6e6c61cc
0340023c
4b40101c
004c111c
06d23664
6d0c70cc
366404c3
00060053
08040c56
ff967016
806c50c3
c037c157
466493cc
746c20c3
0404335c
12c305c3
01963664
08040e56
0336f016
70c3ff96
92c381c3
606c53c3
80378006
20a6cfcc
34c328c3
20c36664
17c4375c
3f866065
61803183
2c6e340b
2c8e342b
2cae344b
0066935c
335c7c6c
07c30404
366412c3
c0760196
08040f56
0336f016
70c3ff96
92c381c3
606c53c3
80378006
20e6cfcc
34c328c3
20c36664
17c4375c
3f866065
61803183
2c6e340b
2c8e342b
2cae344b
0066935c
335c7c6c
07c30404
366412c3
c0760196
08040f56
ff96f016
71c350c3
79ccc06c
2026002c
36644046
326430c3
16546007
0cc7373c
0584255c
235c6d00
4ed20641
60376006
05c39bcc
27c32106
30c34664
0404265c
13c305c3
01962664
08040f56
40c31016
0b08201c
0000211c
6025680c
684c680f
282f63f2
2c2f0053
0b08201c
0000211c
6006284f
700c642f
0361135c
002627d2
1341145c
0872a2bc
724c0133
04c36c0c
0ef4101c
0000111c
08563664
00000804
fe967016
315c51c3
6c0c0644
0010341c
01166af2
0b84301c
0000311c
06c66c0c
80563664
6ccc746c
2006140c
60c33664
335c76ac
255c04c4
2d0017a4
08cb9cbc
2000301c
0800311c
055c7a0f
065c0a01
155c01fd
788017a4
4406788f
600658ce
000678ee
5b8e18af
165c2086
198f01d5
17a4355c
02065980
32c3080d
009e133c
067201c3
1f5c0077
2c0d0021
684d6006
08ad0206
1469155c
19542007
1471355c
01ed365c
1479055c
027d065c
1471155c
32c329ed
049e233c
255c02c3
023c1479
0037302c
00010f5c
01530c0d
301c0116
311c0b84
6c0c0000
366407c6
762c8056
05c38c6c
201c16c3
600600a4
02964664
08040e56
fe967016
606c60c3
000c6ccc
36642006
7aac50c3
04c4335c
17a4265c
9cbc2d00
301c08cb
311c1000
760f0800
178e0506
0a01165c
01fd155c
17a4265c
748f7500
600614ce
000674ee
208614af
01d5155c
365c158f
558017a4
080d0306
133c32c3
01c3009e
00770672
00211f5c
60062c0d
0306684d
165c08ad
20071469
365c1954
69ed1471
033c32c3
10c3049e
1479065c
30ac103c
1f5c2037
2c0d0001
1471265c
01ed255c
1479365c
027d355c
01160153
0b84301c
0000311c
07866c0c
80563664
8c6c7a2c
15c306c3
0148201c
46646006
0e560296
00000804
fe967016
42c360c3
6ccc606c
2006000c
50c33664
335c7aac
265c04c4
2d0017a4
08cb9cbc
1000301c
0800311c
960f43a3
0a01065c
01fd055c
17a4165c
748f7480
54ce4546
74ee6006
14af0006
2086578e
01d5155c
365c158f
558017a4
080d0346
133c32c3
01c3009e
00770672
00211f5c
60062c0d
0286684d
2e0608ad
365c29cd
60071469
065c1954
09ed1471
133c32c3
21c3049e
1479165c
312c213c
2f5c4037
4c0d0001
1471365c
01ed355c
1479065c
027d055c
01160153
0b84301c
0000311c
07466c0c
80563664
8c6c7a2c
15c306c3
01c8201c
46646006
0e560296
00000804
0136f016
50c3ff96
72c341c3
04c4805c
6ccc606c
2006000c
60c33664
335c76ac
255c04c4
2d0017a4
08cb9cbc
311c6006
43a30048
455c9a0f
465c0a01
055c01fd
780017a4
2346788f
400638ce
600658ee
3b8e78af
465c8086
798f01d5
17a4055c
21465800
32c3280d
009e133c
867241c3
0f5c8037
0c0d0001
284d2006
68ad6146
88cd8026
090d1166
04e4355c
28d22c4b
2c3232c3
044e233c
812c213c
055c4c0f
76ac0584
0484335c
2d00588c
00c4301c
48c3640e
60277049
355c0994
6c0c0604
73e427c3
23c30d35
355c0173
602713a1
27c30894
7fff731c
201c0335
442e7fff
844e808b
446e40ab
648e60cb
6c4c762c
16c305c3
01963664
0f568076
00000804
40c31016
06a4305c
1e00233c
6025688c
68cc688f
28af63f2
2c0f0053
600628cf
01e6640f
1341145c
087300bc
145c01e6
a2bc1341
08560872
00000804
60c3f016
f0cc800c
0519105c
402624d2
0515205c
145c184c
2cbc0544
00070880
345c6e94
60070a83
345c6a94
6c6c0604
0014533c
6394a007
08958ebc
08c7045c
0a69145c
341c31c3
60070003
301c1994
311c0448
6c0c2010
0014533c
6dcc70cc
366404c3
1384245c
09c3125c
341c31c3
66d20002
0a24325c
0100331c
70cc2294
06c36d6c
145c3664
31c30a69
0003341c
35946007
03d1365c
13946047
11940007
0624365c
60276e29
345c0c35
60251924
1927345c
04c37c2c
0a61145c
03533664
1489245c
1444145c
245c68a0
282c2524
61476c80
345c0bb4
60251904
1907345c
6d2c70cc
2046100c
70cc3664
04c36d4c
a5d23664
6c6c78cc
366406c3
08958ebc
08e7045c
365c6006
345c0515
001c06c4
011ceb10
2c4c0009
301c4066
311c0fe4
6cac0000
08745abc
08040f56
fd96f016
72c360c3
b80c03c3
7000301c
2010311c
233c4006
401c016f
411c7800
24c32010
f79432e4
725c301c
2010311c
8c0e8a26
8c0e6045
8c0e6045
201c6045
4c0e0090
8f466045
60458c0e
4c0e4c86
15942047
580c75cc
80378026
20772206
02c38d4c
201c17c3
211c7124
69062010
75cc4664
05c36d0c
02f33664
40b74246
7124101c
2010111c
01934006
259d303c
401c640e
842e3f3f
323c2085
23c30010
60972364
f31423e4
72d6301c
2010311c
2c0e2006
2c0e6205
0430301c
2010311c
0332201c
321c4c0f
2c0e6e26
81666045
265c8c0e
321c0923
4c0e0098
0f560396
00000804
61c3f016
201c72c3
211c0c02
501c2010
511c0c04
401c2010
411c0c06
20062010
1c54c007
341c600c
6fd20001
0243305c
305c680e
740e0253
0263305c
303c700e
325c108c
dfe5fff6
41052025
8105a105
043417e4
017c021c
0f56fc93
00000804
0136f016
705c50c3
405c1564
17c308a4
601c4006
611c4000
04c32010
0200431c
001c0335
823c0200
355c180c
83840504
6c2c38c3
c40f642f
787230c3
4025644f
0074323c
7d806412
d800646f
27c9355c
053423e4
22059020
e0948007
200c323c
5d807e05
6e72684c
8076684f
08040f56
40c33016
1564505c
211c4006
680c2010
680f6d92
093124bc
71cc900c
04c36d0c
25c33664
301c2364
311c0098
4c0e2100
808c253c
4c0e6045
311c6946
201c2100
4c0e0085
345c6026
0c5605a7
00000804
800c1016
6cec622c
366404c3
00a8201c
2010211c
6572680c
70cc680f
04c36dac
706c3664
0584335c
366404c3
08040856
40c37016
08a4205c
1564505c
04c4305c
000615c3
c007cc89
001c1094
011c4000
145c2010
b0bc05a4
301c08cb
311c0098
4fe62010
04134c0f
c40c642c
313cc42f
0025087f
27c9345c
f71403e4
236425c3
0098301c
2100311c
253c4c0e
6045808c
69464c0e
2100311c
0085601c
700ccc0e
235c4026
0e5605a7
00000804
0336f016
91c350c3
23642217
036403c3
455cd5ec
323c0644
60070024
700c4d94
0010341c
48546007
0014323c
44946007
303c25f2
60074004
30c32394
2000361c
0b4b333c
233c500c
500f09db
0804323c
32c364f2
700f7972
323c500c
6fd200f4
ed4b61d7
833c37c3
283c208c
500f0a1b
1004323c
32c364d2
700f7972
203c2af2
700c4004
777243d2
323c0073
700f0ddb
79c3782c
0784075c
366414c3
05c3780c
500c3664
200632c3
0010111c
64d23183
749232c3
c076700f
08040f56
3f36f016
60c3e196
43b781c3
ebd76377
05430f5c
cf5c0337
df5c0563
1f5c0583
22f70603
17c4365c
0030233c
a41ca2c3
3a3cfffc
336402c0
986c6577
ba4c8637
180ca677
305c06b7
433c0504
83f70014
2583bf86
610008c3
465c6c10
2bc30644
111c2006
21830010
0564165c
14544007
02b9205c
17c7323c
938491c3
628c09c3
0584165c
7aac4ca0
0464335c
0230141d
a02604f7
91c30093
52c344f7
6c0c798c
0002341c
261768d2
0844315c
18c306c3
366427c3
02c34317
0001041c
27940007
1469365c
23546007
1471165c
17c7313c
0564265c
640c2d00
0001341c
17546007
215c7c0b
41370243
119432e4
215c7c2b
41370253
0b9432e4
315c5c4b
23e40263
365c0694
4ccc2544
4ccf4025
2684265c
6025680c
700c680f
1010341c
1010331c
304b0594
602531c3
0007704e
40062b54
0965265c
341c700c
6ed20010
34c38317
0002341c
a8d269f2
6cac79ac
041c0cc3
16c32000
265c3664
32c30c73
0040341c
e4dc6007
a0070036
0036b2dc
341c3cc3
60074000
59c32254
67327409
1d946007
a0076bf3
06171a94
182c61cc
40c62026
30c33664
60073264
003532dc
31c32317
0002341c
c4dc6007
46570034
06c3684c
2dc318c3
68933664
43c36317
0002441c
800786f7
3c3c2294
60070804
58c31e54
3d8438c3
30c30d8b
000f341c
653703c3
215c19c3
32c30ba3
341c3063
6fd20001
688c4657
155c06c3
82d702b9
241c24c3
36640fff
639304d2
a537a006
03203a3c
65b73364
03f4ab3c
0a24365c
0001341c
5e946007
200b0b97
341c31c3
265c0001
65d22684
602568ac
009368af
6025688c
43d7688f
2b544007
1623465c
341c34c3
60070001
ab972494
10c31409
0001141c
2f5c22b7
2f5c0141
66570005
06c38d8c
459758c3
28c33500
46643ac3
526450c3
e4dca007
786c002d
1663265c
80378206
06c38e0c
00c5101c
466435c3
0007bf5c
a077ab57
00479f5c
81ac0657
18c306c3
3dc34026
40264664
440d2397
60376b97
411c8006
b4830300
0027bf5c
950ca657
18c306c3
23c36317
46643cc3
49c35633
341c700c
60070001
002ab2dc
2684365c
40254c2c
a0264c2f
06d7a5f7
44dc0007
3c3c0029
1c3c0804
60078004
20c31954
46d72dd2
31c32517
49c36685
359d343c
05c3a2d7
029430e4
251745d7
668531c3
49c3a2d7
371d543c
05f70026
46d70253
46d72ad2
315c19c3
82d703c3
35e454c3
45d70294
09c322d7
03c6105c
65f76006
22dc4007
365c0026
4c4c2684
4c4f4025
3cc34cf3
1000341c
57ec59c3
400768d2
32c31974
77ef7f72
01136046
12154007
7f9232c3
6bef29c3
a6576026
06c3946c
125c28c3
a4d702b9
11ac253c
0480393c
1bc34664
011c0006
10830040
20072437
3c3c1654
68d21004
01003d3c
65773364
00a03d3c
3c3c0153
69d22004
00403d3c
65773364
01003d3c
65b73364
fea03d3c
736473c3
20063bc3
0060111c
41c33183
089434e4
0002a21c
fffca41c
77805ac3
04170133
a21c0ad2
a41c0002
1ac3fffc
73c36780
01937364
17c4365c
5f866065
61853283
65773364
336460c5
0bc365b7
511ca006
05830200
05d20477
00e0373c
736473c3
00065bc3
0300011c
2b975083
a0772037
890c4657
18c306c3
23c36317
46643cc3
a0c6a6d2
545c48c3
011302a6
8c2c794c
1bc308c3
36c34357
08c34664
02a3105c
341c31c3
60070004
001a42dc
04042c3c
20544007
325c29c3
602702a1
a6970594
0361555c
3c3ca6f2
60070804
001bf2dc
0007bf5c
00770b57
00479f5c
85ac2657
18c306c3
3dc34006
60264664
680d4397
7aac35b3
0404335c
9f866065
7da03483
58c33364
b580742e
0100373c
d364d3c3
21322557
e132e597
07004f3c
015304c3
03944067
00b317c3
0010313c
136413c3
38c30045
159d333c
323c600e
23c30010
40c72364
0cc3ee94
4000041c
41540007
03832f5c
341c32c3
09c30001
123c400c
63f22a0b
288b123c
17c4365c
5f866065
233c3283
3b3c0200
698003f4
418008c3
00a4313c
28496dd2
280b01c3
402c313c
684b748e
086b74ae
742c14ce
141c0173
742c0001
280b29d2
084b348e
286b14ae
797234ce
313c0073
742f0e5b
265c548b
74ab0766
0776365c
065c14cb
00b30786
303c742c
742f0e5b
17c4365c
3f866065
08c33183
2a8428c3
c35c6980
2d3c015c
323c088c
6180080c
013f143c
016f133c
07c00f3c
41e410c3
48c3f894
02a3045c
341c30c3
60070002
323c4754
343c0060
101c359d
111c8e88
21c30000
105432e4
04a4365c
6cd26c0c
2544365c
40254c8c
66974c8f
0361335c
04dc6007
83d70010
2a548007
1623065c
341c30c3
60070001
2b972394
32c34409
0001341c
4f5c6277
4f5c0121
06570005
06c3818c
659728c3
3ac32980
70c34664
e0077264
000df4dc
265c786c
82061663
8e0c8037
101c06c3
37c300c5
7aac4664
0404335c
1f866065
18c33083
6c80240b
4e204dc3
323c740c
740f601b
08c320a6
0286105c
40a6740c
1b1b323c
740f6f92
542e4006
6ed266d7
0799465c
065c95ed
04b70791
02411f5c
041c35cd
0537000f
48c30273
02b9345c
051775ed
04d710c3
20ac103c
1f5c2237
35cd0101
079d365c
265c55c9
40060795
400c3c3c
4096331c
40260294
323c742c
2b3c0e9b
323c0dcb
44170a1b
323c5632
44570a5b
323c5932
13c30a9b
103c05d7
342f0e1b
451708d2
668532c3
243c49c3
0093359d
205c09c3
443203c3
323c31c3
742f631b
335c7aac
233c0404
7f860030
41f72383
00e14f5c
a205948d
17c4265c
00063bc3
0020011c
60073083
323c1454
3f860030
61853183
698028c3
405c0617
06c30764
4c2b2c0b
03644664
065c140e
00931366
1363165c
4b57340e
542e480b
045c49c3
30c30463
143c6a45
352e359d
27a3265c
365c554e
756e27b3
962d9766
055c58c3
303c02a3
69d20024
20090397
21b72072
00c12f5c
0413400d
0044303c
1c546007
0014303c
18946007
8c096397
541c54c3
a17700fd
00a11f5c
200d0397
461701b3
182c69cc
21c32026
30c33664
60073264
ffd9d4dc
1f96b773
0f56fc76
00000804
3f36f016
60c3f296
42b751c3
024c6277
365c0377
20060664
365c2f8d
133c17c4
5f860030
74801283
0ac34c10
355c1ed2
23c30873
748063d2
323c4c2c
1f86708c
63373083
165c64f2
23370564
42976046
3ac3680d
011c0006
30830010
23176fd2
0564365c
7aac45a0
0444335c
1230141d
2f5c2237
255c0101
2ac302bd
311c6006
23830040
4b544007
00063ac3
0020011c
60073083
365c1a54
606517c4
31833f86
e68b3580
0280233c
936492c3
0240233c
b284b5c3
02c0233c
c284c5c3
75806645
d15c62f7
045301f3
20063ac3
0100111c
60073183
365c1a54
606517c4
32835f86
e50b3580
0100233c
936492c3
00c0233c
b284b5c3
0140233c
c284c5c3
75806345
d15c62f7
00530133
1cc30013
82c3440b
0001841c
265c4006
03b32647
00063ac3
0200011c
60073083
365c1554
606517c4
31833f86
93c36185
c5c39364
393cc984
75800060
72c362f7
801cd2c3
b2c30002
00130053
892c4357
15c306c3
62574297
20c34664
4f940007
0a44365c
11546007
0007af5c
0027bf5c
60b76317
81ac0357
15c306c3
466439c3
22974026
0773440d
0014383c
365c6af2
03c31489
01f70025
00e11f5c
148d165c
00c4373c
05546107
0024383c
12546007
00068f5c
00267f5c
00469f5c
0067bf5c
0087cf5c
617762d7
00c6df5c
80cc0357
8f5c0233
7f5c0006
9f5c0026
bf5c0046
cf5c0067
22d70087
df5c2177
435700c6
06c388ec
429715c3
46646257
fc760e96
08040f56
3f36f016
50c3f996
413761c3
02e4bf5c
02437f5c
02634f5c
02830f5c
855c00f7
55701384
21b7346c
140cb650
17c4355c
5f866065
79803283
3cc38c10
111c2006
31830010
0564155c
265c66d2
323c02b9
258017c7
00c0301c
355c782e
606517c4
32835f86
4e6b7980
7f8532c3
0200331c
001ca5dc
00c4343c
54dc6007
355c001a
60071469
255c2f54
323c1471
93c317c7
0564255c
29c39284
341c680c
60070001
3bc32154
19c34c0b
0243315c
1b9423e4
4c2b3bc3
315c19c3
23e40253
3bc31494
19c34c4b
0263315c
0d9423e4
0014373c
6af2e026
2544355c
40254ccc
e0264ccf
91c30073
343ce006
331c0ff4
14540080
0080331c
680708d4
0010f2dc
94dc6a07
19f30014
00a0331c
001162dc
00c0331c
001404dc
105c2213
27d20cb9
1504355c
40074d09
001704dc
6c0c758c
0001341c
746c68d2
0844335c
16c305c3
36642bc3
045c48c3
30c309c3
0010341c
73546007
17c4355c
0030233c
21833f86
0400323c
80ab1980
341c34c3
60070100
19c36454
02a1315c
09546027
13a1355c
05546027
1469155c
001322f2
2ac37900
018588ac
12c34e6b
40063b05
01774664
00a14f5c
0fe4201c
0000211c
14548007
345c48c3
657209c3
345c6492
000609c6
b4bc28ac
0ac30873
0026814c
40062026
466435c3
04c30653
b4bc28ac
355c0873
1ac304e4
2c29452c
2d09b1c3
75ac013c
266415c3
04e4355c
b2c34c29
323c4d09
a03775ac
0ac38077
03c3800c
21c32146
46646026
0100201c
215c18c3
415c0a27
34c309c3
ffcf341c
315c6872
0ac309c6
05c3618c
36643fe6
e0070006
19c31354
02a1315c
05546027
1469355c
001362f2
455c8006
750c13b6
06c36c2c
25c32026
355c3664
135c1384
31c309c3
0002341c
28c368d2
0a24325c
0400331c
000952dc
0c73155c
341c31c3
64d20010
d2dc0007
e007000b
000894dc
1469255c
54dc4007
1053000b
0504305c
0001341c
d4dc6007
305c000a
67d20cb9
1504355c
80078d09
000a44dc
6c0c758c
0001341c
746c68d2
0844335c
16c305c3
36642bc3
6454e007
305c08c3
331c0a24
5e942000
255c4006
600613b6
0a27305c
17c4355c
9f866065
61853483
01977980
0764405c
2c0b05c3
46644c2b
0686065c
355c08f3
2c091504
255c25f2
400714e1
305c7054
341c0504
60070001
07136a94
0504305c
0001341c
32546007
3054e007
17c4355c
9f866065
65853483
400b1980
0014323c
39c36ef2
648b2e8c
209432e4
64ab402b
1c9423e4
64cb404b
189423e4
155c2106
42061666
61974037
05c38e0c
00c5101c
60064106
01534664
620c0dc3
16c305c3
366424c3
33540027
cf5c0004
45570007
9f5c4077
3dc30047
05c38dac
400616c3
466460d7
81170026
0433100d
1f946087
2684255c
602568cc
305c68cf
233c0504
40070014
343c1494
331c0ff4
0f9400a4
0007cf5c
00770557
1dc320b7
05c385ac
60d716c3
60264664
680d4117
fc760796
08040f56
0136f016
60c3ff96
52c381c3
ebf2e82c
301c0116
311c0b84
6c0c0000
0098001c
80563664
62f2740c
7fe51004
742c740f
742f6c2c
744f62f2
8cac7a4c
17c306c3
00302f3c
466438c3
00192f5c
0014323c
786c65d2
0404335c
323c00f3
67d20024
335c786c
06c305a4
366417c3
66f2742c
165c0086
b8bc1341
01960872
0f568076
00000804
3f36f016
40c3fa96
53c3c2c3
0644b35c
0664235c
a35c40f7
235c1824
323c1471
93c317c7
0564255c
e0069284
d3c36486
1f13d0a4
04c35009
009e303c
813c60b7
38e4ffe0
000f25dc
0010603c
b2dc4547
4547000d
40a707b4
45071054
000df4dc
4ec71b93
000da2dc
00dd231c
000b62dc
44dc45a7
1493000d
20071cc3
000cf2dc
04c4355c
32c34ce9
0001341c
19546007
315c19c3
701202b3
5e7223c3
70801dc3
412c333c
00b8201c
2010211c
455c680f
8ebc06e4
108f0895
06e4355c
2caf2ccc
355c7809
58291336
1323355c
075432e4
1326255c
6c0c760c
366405c3
680c40d7
ffe0101c
0001111c
6af23183
1333255c
49f24037
00011f5c
2dad3ac3
60060093
69ad2ac3
1323155c
402624f2
1326255c
1323255c
1333355c
051432e4
fff0323c
1336355c
0c73255c
341c32c3
6ed20010
08958ebc
15a7055c
355c6006
778c15c7
2c8f2006
2544355c
75cc2ccf
05c36c0c
12e4155c
36644006
1547055c
255c4026
355c0985
6c0c0644
0010341c
56546007
6ccc756c
366405c3
00070077
746c4f94
06c38ecc
00413f5c
39c313c3
02b3235c
466435c3
640c1bc3
323c4057
640f0adb
00213f5c
1525355c
155c0286
a2bc1341
02860872
1341155c
087300bc
1cc305f3
2c942007
201c0116
211c0b84
680c0000
36640886
04538056
101c780c
111c5000
21c302f2
1a9432e4
13c378c9
000f141c
355c2137
31e41499
3f5c1154
355c0081
0173149d
21773809
14a1355c
065431e4
00a13f5c
14a5355c
28c3e026
29a06097
20279980
fff085dc
069607c3
0f56fc76
00000804
03c3600c
0524135c
1000233c
08f118bc
00000804
0136f016
105cfe96
a00606a4
65c375c3
100c273c
6d0063ec
6006656f
01b36037
83ac63ec
e0258d61
6a0563ac
601763af
802543c3
40858037
0141315c
84c38017
ef1483e4
00012f5c
014d215c
100c463c
0404305c
658f6e00
60776006
305c0293
43cc0404
c0254e61
63cc02b0
225c28c3
6d000684
605763cf
821c83c3
8f5c0001
80850027
0151315c
82c34057
e81483e4
00212f5c
015d215c
a025a5af
0354a187
f6f32785
80760296
08040f56
0136f016
73c362c3
41c30364
a80c4364
81c32c0c
25c30212
00d334c3
027f213c
7fe54800
7bf23364
428d303c
780f7580
100c343c
698028c3
80767c0f
08040f56
02c330c3
480c1364
2c6e4c0f
313c2c4e
6980100c
0804600f
40c37016
0644005c
16e4645c
145cb06c
313c1471
145c17c7
4c800564
341c680c
60070001
345c1d54
60071469
125c1954
200702a1
400c1594
341c32c3
66d28000
6e7232c3
0bdb313c
355c600f
04c307c4
38093664
355c25d2
04c307a4
716c3664
04c36c4c
0e563664
00000804
40c33016
1384205c
09c3025c
341c30c3
66d20002
0a24325c
0100331c
345c3994
64f213c3
13e7345c
8ebc0673
50c30895
13e4145c
045c24f2
055313e7
0ad3245c
0014323c
323c65d2
60070024
54a02194
13c3045c
001c10c3
011c4240
313c000f
23e4028d
706c1535
102c6dcc
40862006
30c33664
6cd23264
13e7545c
0904345c
345c6025
722c0907
04c36f6c
0c563664
00000804
3f36f016
60c3fd96
d1c372c3
8870d264
16e4825c
1353925c
17c4325c
3f866065
68053183
a384a0c3
60073dc3
0008f2dc
408b0ac3
375c4a12
32e412e4
275c1254
7e0c12e7
07c36c0c
375c3664
4c091504
3ac348f2
301c4c8b
311c08c4
4c0f2010
1471075c
17c7303c
0564175c
375cac80
606517c4
32835f86
79806185
405c0cc3
07c30764
4c2b2c0b
03644664
04f6055c
32c357ec
111c2006
31831000
32c36ad2
77ef7c92
0bb6055c
255c4006
01330bc6
0bb3155c
0037313c
62526180
0bb6355c
682b28c3
333c67d2
61800037
682e6252
38c30073
931c0c2e
0f5400ff
0bb3255c
0bc3155c
608009c3
05d423e4
610009c3
031531e4
0bc6255c
0784865c
0863565c
bf3c7e2c
8cec00a0
265c05c3
365c0873
29a00743
3bc34006
90c34664
7e2c9364
05c38cec
21c32006
46643bc3
2ac30364
482c680c
20372026
1cc3e077
0784415c
042019c3
38c313c3
5d0c4664
17c4375c
1f866065
79803083
0a3c880c
4e6b00c0
3b0512c3
37c32dc3
03964664
0f56fc76
00000804
50c33016
8ebc41c3
145c0895
40a015e4
15e7045c
0ba4145c
345c6880
32e40ba7
345c0634
60250bc4
0bc7345c
0ba4345c
145c740f
342f0bc4
08040c56
41c37016
c15752c3
0b67165c
0b87265c
08cc201c
2010211c
4085280c
65a0480c
33646180
34e46e00
a0250234
0ba7365c
0bc7565c
08958ebc
15e7065c
08040e56
336430c3
716c201c
2010211c
301c680e
311c8004
2c0b2010
241c21c3
0047f9ff
00870854
00270854
251c0794
00930600
00534a72
301c4972
311c8004
4c0e2010
00000804
0ae4305c
305c31a3
aabc0ae7
08040904
0736f016
91c370c3
335c600c
a3c30361
21546007
2fc30416
a2c34085
513c2056
8e24ffc0
0086f524
08cc78bc
04a4355c
0400441c
60066bd2
04a7355c
82bc0086
800708cc
f3242754
008604b3
08cc82bc
f32482d2
0080693c
853ca026
383c0014
163c0010
2dd23a1d
8d0c7c6c
400607c3
46643ac3
62d238c3
a025c185
ee94a0c7
2c6c39c3
7c6c27d2
07c38d0c
3ac34006
e0764664
08040f56
3f36f016
d0c3f896
c2c351c3
005c6037
00770444
20b7258c
4137562c
341c32c3
331c0580
07540180
0400331c
331c0454
21940100
6972760c
2117760f
241c21c3
301c000f
311cc750
233c0011
41b72a1d
4000231c
101c0435
21b74000
32c34097
0098321c
73c361f7
8006a177
b4c364c3
0833a4c3
0263155c
000b0cc3
233c6420
0cc3fff4
23e4606b
0cc37c15
091944bc
c0268006
0f73b4c3
233c38c4
393c0034
a2c3100c
8f5ca384
c00700e4
853c2254
2dc30540
8d8c6a2c
15c30dc3
0040253c
466438c3
235c6157
355c01f1
23e401f1
760c7194
111c2006
31834000
6a546007
235c6157
355c01e9
23e401e9
a1776394
78c347c3
0263155c
2cc320f7
6520480b
fff4233c
606b0cc3
3a1523e4
32c35c6b
1fff341c
0040933c
3dc389c3
0303035c
838430c3
3bc3c8d2
38843a84
21c32197
2d1423e4
03c36057
225460e4
3a843bc3
b884b3c3
20170dc3
39c34117
091a7ebc
0cc390c3
13c360d7
091944bc
373cc6d2
702e108c
100e0026
108c293c
323c7c2c
7c2f3a1b
b40cc025
8f94a007
c7f247c3
20974006
0636215c
02d3a006
b35c6097
635c0626
c0270636
702c0554
702f6f72
20970173
04e4315c
0bdb363c
04e7315c
47c30073
05c3fd93
fc760896
08040f56
fe96f016
505c40c3
c1cc1824
205c4006
606c1887
0524335c
14c30fc3
740c3664
0d204017
09740007
47d25589
23c3744c
073502e4
758d6006
04c378cc
36641fc3
045c03f2
029612e4
08040f56
30c3f016
505c41c3
205c0644
000c0664
635c204c
315c0544
60470161
80260294
341c7869
68f20001
205c4026
61cc0ab5
36646dcc
800704b3
680c1494
0001341c
1e546007
6007684c
682c1b94
711ce006
37830001
740c66f2
000f341c
10546007
2006740c
0060111c
40063183
0040211c
37e472c3
622c0594
6cac3809
0f563664
00000804
0361205c
62cc45d2
6c0c6c0c
08043664
0136f016
08c8301c
2010311c
305c8c0c
4c291504
0604305c
341c6c6c
66d20010
305c44f2
23c31771
605c5fe5
701c0584
711c08c4
00932010
500c353c
323c9180
79800cc7
0641135c
bc0c2cf2
305c4025
83c31771
ffff821c
ef3528e4
fdb321c3
807604c3
08040f56
0736f016
40c3ff96
13c361c3
736472c3
62ac3890
0484335c
40b0731c
59090894
008502c3
2f5c0037
590d0001
4c0009c3
2af201c3
01e9165c
17c7313c
0564045c
033c6c00
165c0480
313c01e9
83c317c7
0564145c
38c38184
345cae8c
6c0c0644
0104133c
1000301c
31c322f2
680e37a3
284e200b
a21ca0c3
3ac30002
686e6c0b
133c30c3
288e023e
28ae348b
28ce34ab
28ee34cb
00a4731c
200b1c54
0ac3290e
092e000b
294e2c0b
16c4345c
696e6412
341c7a0c
65d21000
61c909c3
698e6432
282e2006
16c4345c
345c6025
013316c7
105c08c3
31c302b3
c000001c
682e30a3
6c8c722c
16c304c3
01963664
0f56e076
00000804
40c31016
0b1c201c
0000211c
6025680c
684c680f
282f63f2
2c0f0053
0b1c301c
0000311c
60062c4f
03c3640f
1341145c
0872a2bc
08040856
60c3f016
52c341c3
0e26e00c
08cc78bc
542c702c
704c64d2
00534c2f
544c502f
700c504f
6d00540c
6006700f
744f742f
0e26740f
08cc82bc
00467c4c
301c2c0c
311c0fe4
4d0c0000
08c8d4bc
165c0026
b8bc1341
786c0872
06c36e6c
0f563664
00000804
000c1016
0544305c
4c29208c
8f4c4612
335c6a00
60870424
640c0394
61070093
642c0494
01533664
301c0116
311c0b84
6c0c0000
366406a6
08568056
00000804
0336f016
50c3fe96
40372077
e00c93c3
6ccc606c
202607c3
40c33664
000780c3
80c35354
17c4355c
0030133c
12835f86
375cc080
63d20361
08cb9cbc
06c37eec
9cbc2f0c
904f08cb
01231f5c
355c56ac
606517c4
30831f86
04a4025c
65806c00
56ac70ce
17c4355c
1f866065
025c3083
6c0004a4
700e6580
17c4355c
5f866065
702e3283
345c6026
00860296
0286045c
313c780c
4086601b
231b323c
2f5c780f
584d0021
6bf26057
60877f2c
275c0894
45f20361
0724375c
784f6105
0066965c
00013f5c
08c379ed
c0760296
08040f56
00000034
00000038
0000003c
00000040
00000064
00000068
0000006c
00000070
00000074
00000078
0000007c
00000080
00000084
00000088
0000008c
00000090
01000001
03030202
226420c3
011c0086
200b2200
1000301c
31a33223
600e3364
00000804
606cfb96
6ca0204c
141d404b
20b71320
00413f5c
1f5c60f7
202d0061
03356507
602d6506
01732006
61004117
00811f5c
0185135c
40774025
00211f5c
60292137
12c34117
f1b431e4
7fe532c3
1f5c6037
200d0001
08040596
60c37016
26f251c3
0004f524
00040004
872b0013
fff0343c
436443c3
243c798c
6c2c0010
153c06c3
36642e1d
0e5694f2
00000804
0136f016
26f270c3
0004f524
00040004
513c0013
244f0040
83c36e24
8006f524
0014643c
0010363c
3a1d153c
7d8c2ad2
07c36c2c
c2d23664
8025a185
f19480c7
4004383c
f32462d2
0f568076
00000804
40061364
31e46009
40260214
080402c3
0736f016
70c3fc96
82c3a1c3
20d08364
680929c3
6c546007
7fe5484b
228d333c
667438e4
19c348c3
68a02469
83e47e05
43c30235
7d8c4364
00c05f3c
07c36c0c
366415c3
d84fc0d7
2c697ccc
620531c3
78ce7180
6c697ccc
2ac3782e
865cc80f
18c30006
43c36620
801c4364
07530001
6c0c7d8c
15c307c3
383c3664
40d70010
3f9d263c
0c4b39c3
24c314c3
30c32364
23e43364
10c30235
236421c3
180c383c
4cce7980
0010383c
363c6077
60073e1d
56c31294
017343c3
6c2c7d8c
340c07c3
243c3664
40370010
00014f5c
48e4a105
01d3f414
00211f5c
826481c3
43c37120
80074364
865cc694
80b70196
40260073
3f5c40b7
03c30041
e0760496
08040f56
ff96f016
61c340c3
72c36364
53c37364
618c5364
1fc36c0c
40173664
0c6970cc
484f2800
0c6970cc
620530c3
68ce7580
0c6970cc
620530c3
680e7580
6c6970cc
6026682e
00c66b2e
c4ee0b0e
551ce42e
a40e6000
019602c3
08040f56
60c37016
968ca14c
30c34664
063c544c
13c30500
0e562664
00000804
22641364
0cac600c
0f944027
00ff131c
40060594
0996205c
323c0213
33e3100d
0993205c
00f33283
602648f2
205c3123
32a30993
0996305c
00000804
400e4006
202e2026
4106404e
101c406e
204f03e8
00000804
301c3016
311c01e4
8c0c4102
434c9ff2
60262a4c
3523a009
318333e3
301c6a4f
311c01e4
8c0f4102
08040c56
60a04006
027432e4
02c34026
00000804
080400a0
40c31016
78bc0f26
334c08cc
6026464c
30231009
664f32a3
82bc0f26
085608cc
00000804
ff96f016
62c351c3
103c83c6
03130040
4007440c
742c0815
640f3203
f40c600c
600f3703
233c640c
440f080c
6007600c
32c30415
640f6072
6112600c
343c600f
6037fff0
00014f5c
00ff431c
402ce294
600c582f
0196780f
08040f56
fa963016
101c51c3
111c54fc
340fbbcc
201c45c3
211c8d96
243c8384
600c027e
001c23c3
011cffff
208300ff
3da9101c
8571111c
00a620b7
200600f7
0080111c
12c33183
011c0006
10032c00
12c366d2
311c6006
13031300
323c500c
1303108c
100c313c
00066177
23030137
6097500f
188c233c
333c60d7
60f7e92c
111c2006
20b72000
01000f3c
00801f3c
d2bc2fc3
20570941
7e326017
11ac213c
3203740c
313c740f
500cf08c
700f3203
0c560696
00000804
31c3ff96
60e73264
7f851335
01732180
640c400c
088d223c
088d333c
027f303c
fe7f213c
0030303c
f3b413e4
7fe501b3
01532180
60376009
203c4409
3f5c00df
313c0001
01e4ffdf
0196f614
00000804
240c31c3
2c4b200f
0804204e
ff961016
4026600c
840c4037
32e424c3
60060994
404b6037
23e4644b
20260354
2f5c2037
02c30001
08560196
00000804
50c37016
000641c3
019310c3
188c213c
0074313c
363cd522
341c308d
01800001
14e42025
0e56f414
00000804
31c3ff96
60373264
600648d2
00011f5c
602521a1
fb9423e4
08040196
47d21016
85a26006
602581a1
5cf25fe5
08040856
f5244e24
69d2600c
7fe5600c
602c600f
602f6c2c
604f62f2
4004323c
f32462d2
00000804
f5244e24
6025600c
604c600f
202f63f2
2c0f0053
6006204f
323c640f
62d24004
0804f324
f5244e24
68d2600c
600f7fe5
6c0c602c
62f2602f
323c604f
62d24004
0804f324
f5244e24
6025600c
604c600f
202f65f2
640f204f
602c0093
202f640f
4004323c
f32462d2
00000804
8e243016
600cf524
14546007
600f7fe5
4006602c
23c30073
13e46c0c
46f2fd94
4004343c
f3246bd2
240c0133
404f22f2
343c280f
62d24004
0c56f324
00000804
40c37016
ce2451c3
0ce6f524
08cc78bc
6025700c
704c700f
b02f63f2
ac2f0053
6006b04f
0ce6742f
08cc82bc
4004363c
f32462d2
08040e56
fa961016
326431c3
22646177
412c4137
215768a9
43c327d2
80f78072
00611f5c
43c300d3
80b78092
00411f5c
68a928ad
88d28117
217213c3
3f5c2077
68ad0021
43c300f3
80378192
00011f5c
616c28ad
6c0c406c
0110023c
00a12f5c
4f5c12c3
24c30081
06963664
08040856
32c3fd96
32641364
0a946047
313c402c
294c01c7
6c8c6c80
0348335c
5fe602b3
602740b7
400c1e94
0487313c
6c80282c
2c286c8c
60e8022c
081513e4
207725a0
00213f5c
60b73064
01080193
40b74006
07f410e4
20372420
00011f5c
20b71064
00412f5c
039602c3
00000804
31c3fc96
22643264
67d22009
617231c3
3f5c60f7
00d30061
619231c3
3f5c60b7
600d0041
47d22009
627231c3
3f5c6077
00d30021
629231c3
3f5c6037
600d0001
08040496
c0967016
536451c3
6c09612c
2006406c
00051f5c
4f5c89e9
1fc3000d
c42eca6b
0014433c
600c85d2
cc296c8c
602c0093
cd896d2c
00256f5c
315c6a2b
88d2002e
6c8c600c
10f3435c
003e415c
602c00d3
cf6b6d2c
003e615c
8c6c614c
2fc315c3
46646126
0e564096
00000804
bf967016
612c1364
806c6c09
10402f3c
523ca006
d28b805e
000e625c
0014633c
c7d2c037
6c8c600c
5f5cade9
00b3003d
00016f5c
003d6f5c
684e7209
686e7209
8c6c614c
00402f3c
46646106
0e564196
00000804
0736f016
50c3c096
a1c382c3
804ca364
612c2250
063ccc09
10c30014
740c03d2
763c2c0c
67c30024
742ce3d2
28c3cc0c
700e6869
23c36889
38c3702e
704f6ca9
444d0bd2
454e506b
658e706b
68ec29c3
084c6d0c
edd23664
784d7049
594e506b
798e706b
68ec29c3
084c6d0c
366416c3
10003f3c
233c4006
554c805e
05c3886c
2fc31ac3
46646026
e0764096
08040f56
40c33016
618c51c3
36646c0c
6c4f740c
486950cc
20e64c2e
40262f0e
233c4f2e
70cc0100
08802c69
08040c56
13647016
3ff4513c
6c6961ec
051435e4
333c61cc
00735a1d
6cac614c
0e563664
00000804
c0963016
3f3ca026
533c1000
414c805e
2fc3886c
466435c3
0c564096
00000804
40c3f016
136462c3
3ff4513c
6d8b620c
0c3535e4
ec09612c
341c37c3
66d20002
6c2c602c
5a1d333c
714c00b3
04c36cac
366426c3
08040f56
0336f016
40c3ff96
612c81c3
414cec09
60aca44c
10c30d09
20372025
00010f5c
153c0d0d
013c083e
673c508c
cdd20014
6cac700c
0969335c
07946027
36940067
3ff4313c
32946067
1b540087
08b40087
11540047
13b40047
24940027
00c70153
00c71454
01071014
07e71354
02b31b94
0333696c
1654c007
02b3698c
027369ac
023369cc
01f369ec
6a0ccdd2
373c0193
68d20024
00f36a2c
04c36a4c
366418c3
68ac00b3
25c304c3
718c3664
04c36c4c
366418c3
c0760196
08040f56
40c37016
612c414c
644cac09
60676dc9
60672f54
602706b4
60470a54
03934494
3f546207
00ff331c
06133e94
366468cc
0014353c
700c66d2
680c4e2c
680f6025
0024353c
2f546007
4e4c702c
31c3292b
692e6025
68ec0513
353c3664
60070014
700c2254
682c4e2c
682f6025
353c0393
69d20014
3664690c
4e2c700c
6025686c
0233686f
6c4c618c
692c01b3
353c3664
69d20014
4e2c700c
6025688c
0073688f
3664694c
08040e56
c0967016
61c340c3
00ac6364
0030123c
b0bc4106
2f3c08cb
60061000
805e323c
ac6c714c
16c304c3
60262fc3
40965664
08040e56
c096f016
71c350c3
4f3c7364
60061000
805e343c
0f3c606c
133c0010
41060060
08cbb0bc
cc6c754c
17c305c3
61262fc3
40966664
08040f56
c096f016
71c350c3
4f3c7364
60061000
805e343c
0f3c60ac
133c0010
480600f0
08cbb0bc
cc6c754c
17c305c3
68262fc3
40966664
08040f56
c096f016
71c350c3
606c7364
10004f3c
243c4006
0f3c805e
13c30010
094282bc
cc6c754c
17c305c3
60e62fc3
40966664
08040f56
bf967016
61c350c3
48696364
206c4037
2f5c4006
3f5c0025
3f5c0001
612c002d
32c34c09
0001341c
600c67d2
4c096c8c
00352f5c
60260093
00353f5c
45f24017
00700f3c
011320c5
23c36017
08944027
00700f3c
41062225
08cbb0bc
0f3c0173
60170070
232523c3
f6544047
9cbc2106
754c08cb
05c38c6c
2f3c16c3
61660040
41964664
08040e56
60c37016
13c351c3
036402c3
75cc1264
ff00433c
23c372a0
542e2364
0100303c
740e6980
03942027
00536046
70ee6066
01e5355c
7000051c
8e24100e
794cf524
063c6c4c
15c30500
343c3664
62d24004
0e56f324
00000804
40c37016
642b2364
af00c44c
cc6970cc
620536c3
64ce6980
cc6970cc
620536c3
640e6980
74ee6086
615cc086
251c01e5
540e7000
f524ae24
6c4c714c
0500043c
353c3664
62d24004
0e56f324
00000804
40c37016
642b2364
af00c44c
cc6970cc
620536c3
64ce6980
cc6970cc
620536c3
640e6980
00ff301c
251c74ee
540e7000
f524ae24
6c4c714c
0500043c
353c3664
62d24004
0e56f324
00000804
fd963016
51c340c3
22645364
32644077
60ac6037
32c34c09
0010341c
19546007
6e6c614c
00801f3c
36645fe6
400d40a6
00212f5c
505c404d
2f5c001e
40ad0001
402d4086
6c0c714c
209704c3
366440c6
0c560396
00000804
fd963016
51c340c3
22645364
32644077
60ac6037
60076c08
614c1915
1f3c6e6c
5fe60080
41063664
2f5c400d
404d0021
001e505c
00012f5c
408640ad
714c402d
04c36c0c
40c62097
03963664
08040c56
fe96f016
51c340c3
72c35364
32647364
353c6037
633c0a0b
60ac0010
31c32c29
0008341c
30546007
6e6c614c
00401f3c
36645fe6
400d4186
00013f5c
505c604d
c047001e
502c0a94
01c7373c
6c80294c
235c6c8c
01330371
373c500c
282c0487
6c2c6c80
0199235c
135c40ad
206e0353
0363235c
6106408e
714c602d
04c36c0c
41462057
02963664
08040f56
fe963016
32c340c3
536451c3
60373264
6ca860ac
16156007
6e6c614c
00401f3c
36645fe6
400d4606
00012f5c
505c404d
4066001e
714c402d
04c36c0c
40a62057
02963664
08040c56
fd96f016
62c350c3
71c343c3
42647364
6e6c614c
00801f3c
36645fe6
200d21e6
0030143c
3f5c2077
602d0021
204d3809
2d0974ac
e04e206d
4d0974ac
3fe512c3
2f5c2037
4d0d0001
6c0c754c
209705c3
366440c6
0f560396
00000804
60c37016
036402c3
880945cc
02548027
a40b8046
7fe535c3
536453c3
203c32c3
243cfff4
233c612c
ac2efeee
7fa565cc
794c65cf
06c38c2c
0040253c
46646026
08040e56
ff963016
51c340c3
614c5364
1fc36e6c
36645fe6
400d4ae6
4046a02e
714c402d
04c36c0c
40862017
01963664
08040c56
fd96f016
72c350c3
61c343c3
42646364
6e6c614c
00801f3c
36645fe6
200d21c6
0030143c
2f5c2077
402d0021
204d2026
001e605c
17c300a5
b0bc24c3
74ac08cb
12c34d09
20373fe5
00012f5c
754c4d0d
05c36c0c
243c2097
36640050
0f560396
00000804
0336f016
80c3fe96
036401c3
40372264
936493c3
1004193c
44542007
4c2c38c3
01c7303c
ac80294c
47c3e006
08c3c046
00401f3c
88bc5fe6
42660944
6026400d
905c604d
4e24001e
c027f524
60171594
202713c3
73290794
002e305c
732d6006
20170293
11942007
305c7349
3f5c002e
734d0001
748c0153
02f9335c
002e305c
2006748c
02fd135c
4004323c
f32462d2
402d40a6
1094c027
4c4c7e2c
4c4f4025
28c30173
303ce80c
5c2c0487
8c4c6d00
c02651c3
18c3f7b3
6c0c654c
205708c3
366440e6
c0760296
08040f56
313c20c3
6412fff0
00066180
001c0c6f
011c0180
0c2fc107
200c313c
01334980
ffe7225c
0180301c
c107311c
ffa7325c
5e053fe5
080436f2
313c20c3
6412fff0
00066180
001c0c6f
011c0180
0c0fc107
200c313c
01334980
ffe7225c
0180301c
c107311c
ff87325c
5e053fe5
080436f2
311c6186
201c4107
4c0e0080
00000804
009c301c
4107311c
0080201c
08044c0e
41866206
4107211c
221c680e
680e0090
00000804
fe96f016
03c340c3
51c3c1d7
300c5364
62056880
f04b602f
7e2537c3
101c6d20
111c7ffe
31839fff
8000201c
6000211c
604f32a3
03932026
200c313c
313c4180
7180180c
e82fec0c
37c3ec4b
701c6025
711c7ffe
37839fff
8000701c
6000711c
684f37a3
0010313c
1f5c6037
16e40001
31c30534
35e43364
313ce014
7e05200c
684c4180
6000351c
67c6684f
2100311c
133c6c0b
60860014
20076077
20c31394
301c2364
311c0092
4c0e2100
808c203c
4c0e6045
311c6746
701c2100
ec0e0085
1f5c2077
01c30021
0f560296
00000804
13641016
0010313c
fffe201c
0001211c
41803283
0180401c
4107411c
111c2606
01134107
700e600b
341c640b
7df20008
02e40045
0856f894
00000804
6746ff96
2100311c
23644c0b
4c0e4672
211c47c6
27c62100
2100111c
341c680b
7ad20040
341c680b
76f20001
233c640b
60260014
4cf26037
311c6406
6c0b4080
0008341c
64d26037
640e6086
3f5c4037
03c30001
08040196
6746ff96
2100311c
23644c0b
4c0e4672
211c47c6
680b2100
0040341c
680b7dd2
0001341c
67c679f2
2100311c
303c0c0b
60370014
00012f5c
019602c3
00000804
ff967016
10c341c3
22641264
311c6006
00064140
0010011c
60060c0f
4108311c
013c4c0e
4006088c
511ca086
01334108
343c740b
623c271d
c0370010
00012f5c
f71420e4
0014313c
608668d2
4108311c
70804c0b
fffd235c
311c6006
c0064108
6086cc0e
4140311c
011c0006
0c0f0010
0e560196
00000804
80c8301c
4103311c
201c6c0b
211c80f4
080b4103
03ff341c
81ac003c
00000804
0d09612c
211c4246
61002040
080c033c
6026400b
100d133c
31c312a3
600e3364
00000804
0d09612c
211c4246
61002040
080c033c
3364600b
123c4026
21e3100d
600e3283
00000804
326430c3
211c4046
680e4107
0804080b
036421c3
301c2264
311c013e
101c4107
2c0e00ff
013c301c
4107311c
61c54c0e
08040c0e
226420c3
311c6006
6c0b4107
141c13c3
6306ffcf
4107311c
0230001c
49f20c0e
201c6045
4c0e0220
02066045
05330c0e
0c944027
311c6346
001c4107
0c0e0210
44066045
24724c0e
40470393
63460c94
4107311c
0c0e0606
201c6045
4c0e0200
01f32572
0d944067
311c6346
001c4107
0c0e0230
00ca321c
4c0e4026
0030151c
311c6006
2c0e4107
00000804
226420c3
013e301c
4107311c
00ff101c
301c2c0e
311c013c
4c0e4107
6c0b6505
201c3364
211c0166
080b4107
81ac003c
00000804
226420c3
013e301c
4107311c
00ff101c
301c2c0e
311c013c
4c0e4107
6c0b6585
080403c3
226420c3
013e301c
4107311c
00ff101c
301c2c0e
311c013c
4c0e4107
6c0b65c5
080403c3
226420c3
013e301c
4107311c
00ff001c
301c0c0e
311c013c
4c0e4107
236421c3
4c0e6105
808c213c
0142301c
4107311c
08044c0e
226420c3
301c1364
311c013e
001c4107
0c0e00ff
013c301c
4107311c
21c34c0e
61454b72
08044c0e
30c3ff96
60373264
60271264
26d21494
00010f5c
013d025c
201c0433
211c8222
680b4103
ff7d341c
4e05680e
341c680b
0273ffef
600625d2
013d325c
201c01f3
211c8222
680b4103
351c3364
680e0082
680b4e05
64723364
0196680e
00000804
12640264
61862df2
4107311c
4c0e4806
211c4006
680b4107
fffe341c
202705b3
61860e94
4107311c
0200201c
40064c0e
4107211c
341c680b
03d3fffd
0e942047
311c6186
201c4107
4c0e0400
211c4006
680b4107
fffb341c
206701f3
61860e94
4107311c
8000201c
40064c0e
4107211c
341c680b
680efff7
013e301c
4107311c
00ff201c
301c4c0e
311c013c
2c0e4107
638509f2
101c4c0b
21a38000
4c0e2364
00270173
201c0994
211c0158
680b4107
7fff341c
0804680e
326430c3
301c6ef2
311c009c
48064107
40064c0e
4107211c
3364680b
06136072
0f946027
009c301c
4107311c
0200201c
40064c0e
4107211c
3364680b
04136172
0f946047
009c301c
4107311c
0400201c
40064c0e
4107211c
3364680b
02136272
0f946067
009c301c
4107311c
8000201c
40064c0e
4107211c
3364680b
680e6372
00000804
10c321c3
22641264
013e301c
4107311c
00ff001c
301c0c0e
311c013c
4c0e4107
6b862af2
4107311c
0096201c
321c4c0e
019300fe
20276006
6b860994
4107311c
0108201c
321c4c0e
001c00fc
0c0e8000
00000804
036421c3
301c2264
311c013e
101c4107
2c0e00ff
013c301c
4107311c
61854c0e
20c30c0e
301c4b72
311c0146
4c0e4107
00000804
226420c3
311c6306
3fe64107
60452c0e
321c2c0e
2c0e0080
2c0e6045
311c6446
25064107
61862c0e
4107311c
1088101c
40272c0e
301c1194
311c00a0
3fe64107
60852c0e
301c2c0e
311c009e
45264107
60854c0e
404701d3
301c0d94
311c00a8
3fe64107
301c2c0e
311c00a6
45264107
08044c0e
326431c3
0e946027
4d8b303c
201c6212
211c4000
6d004114
ffff201c
003f211c
303c01b3
6212450b
4000201c
4114211c
201c6d00
211cffff
0283000f
08040c0f
600cff96
0d947fe7
400f4006
133c30c3
21c3021e
40374025
00011f5c
00732c0d
600f6025
08040196
00ba201c
4107211c
341c680b
65d22000
341c680b
680edfff
010c201c
4107211c
3364680b
680e6872
341c680b
680efeff
00ba201c
4107211c
3364680b
680e6472
00000804
001c20c3
011c010c
600b4107
62723364
280b600e
00fc301c
4107311c
282b2c0e
2c0e6045
6045284b
286b2c0e
2c0e6045
6045288b
28ab2c0e
2c0e6045
604528cb
48eb2c0e
4c0e6045
341c600b
7df20004
00000804
326431c3
6027400b
301c0e94
311c9898
4c0e4103
6045402b
404b4c0e
4c0e6045
00f3406b
989c301c
4103311c
402b4c0e
4c0e6045
9884301c
4103311c
23644c0b
4c0e4472
00000804
ff96f016
61ec50c3
cc4be1ac
00370c49
211c4446
21064107
2186280e
4107111c
840e8106
30c30c8b
0004341c
620666d2
8046680e
0073840e
080e0206
0948b6bc
0948aebc
0014363c
740c69d2
9c0c6c4c
200605c3
01c9235c
363c4664
68d20024
05c37c0c
4f5c2006
24c30001
01963664
08040f56
0136f016
81c340c3
cc8b61ec
a1ace12c
009a301c
4107311c
4c0e4406
2006740c
366421c3
04c3740c
40262006
740c3664
200604c3
36644046
04c3740c
40662006
aebc3664
163c0948
21c3088b
0014363c
313c65d2
23c3f005
363c2364
62d20024
1c094d72
341c30c3
65d20001
62077cc9
43720294
0065323c
00ba201c
4107211c
363c680e
6ad20084
301c5d0b
311c00f4
4c0e4107
60855d2b
64464c0e
4107311c
4c0e4106
311c6186
4c0e4107
648529d2
0610001c
321c0c0e
0c0e0086
660600f3
4107311c
0410201c
61864c0e
4107311c
1000001c
18c30c0e
313c1364
23c3fff0
62062364
4107311c
66464c0e
4040311c
60452c0e
4c0e4006
311c6486
001c4107
0c0e0c35
211c4306
680b4105
62723364
6306680e
4107311c
4c0e5fe6
00c8321c
301c4c0e
311c009e
08064107
60850c0e
60850c0e
62c50c0e
201c0c0e
211c800a
680b4103
63723364
301c680e
311c00aa
40464107
60454c0e
60454c0e
65c54c0e
80764c0e
08040f56
fe967016
536451c3
253c602c
2d4c01c7
580cc880
40774aa9
4af26c6c
00212f5c
00052f5c
21c68cec
605725c3
20060113
00051f5c
21068cec
600625c3
788c4664
0464235c
235c4072
02960467
08040e56
ff961016
236421c3
323c802c
314c01c7
2c8c6c80
0464315c
315c6172
706c0467
1f5c2006
8cec0005
60062186
01964664
08040856
50c33016
618c41c3
36646c0c
6c4f700c
2c6f2006
0140233c
2c6b74cc
0c560880
00000804
fc967016
536451c3
353c202c
454c01c7
4c8c6d00
0444325c
0044633c
68ccc0f7
1254c007
0251235c
40b74172
00414f5c
0255435c
c006646c
00056f5c
21468cec
600625c3
235c0253
40720251
4f5c4077
435c0021
646c0255
00616f5c
00056f5c
20668cec
60d725c3
04964664
08040e56
0136f016
80c3ff96
61c342c3
42646364
363c402c
294c01c7
ac8c6c80
e86c74cc
8027484c
88cc1694
0300033c
0200133c
0080233c
46646305
0464355c
355c6072
60060467
00053f5c
08c39cec
00d320a6
1f5c20c6
9cec0005
26c321a6
46646006
80760196
08040f56
40c31016
336401c3
31a12509
33646025
31c1206b
33646045
31c1200b
33646045
31c1202b
13c36045
604b1364
70c16332
0020313c
51c13364
0020033c
08040856
ff963016
402c51c3
313c24eb
294c01c7
8c8c6c80
6c0c302c
60276ea9
620c1594
245c0ceb
61000393
236423c3
03a6245c
140c9489
74bc34c3
0364094e
80379000
00013f5c
0196748d
08040c56
fe963016
04eb402c
01c7303c
6e80a94c
040c4c8c
6c0c8489
a0066ea9
6027a077
6a6c1a94
000f305c
0281525c
525ca0ad
35c30393
336460e5
0386325c
343c606e
60370070
00015f5c
325ca077
61720404
0407325c
00210f5c
0296048d
08040c56
fe963016
402c41c3
313c24eb
294c01c7
688c4c80
100c2ccc
680cb089
40774006
40074ea9
648c1094
000f305c
205c44ac
64ec002f
004f305c
00c0253c
3f5c4037
60770001
00211f5c
0296308d
08040c56
ff961016
202c21c3
303c08eb
054c01c7
8c8c6c00
2989680c
68892c2d
002503c3
1f5c0037
288d0001
245c4026
700c02e5
7100001c
0002011c
123c4c0b
5cbc0057
045c0a7c
345c0427
6d720404
0407345c
08560196
00000804
0336f016
60c3fe96
402c81c3
303c04eb
294c01c7
ec8c6c80
28c39ccc
925ca80c
6c0c0021
00066ea9
60270077
500c3e94
000f255c
355c702c
045c002f
055c0263
79ac004e
01066c2c
0080143c
36644046
6c2c79ac
143c0086
40460180
304c3664
005f155c
255c506c
70cc007f
009f355c
0160193c
2f5c2037
40770001
001c7c0c
011c7100
4c0b0002
0057123c
0a7c5cbc
0427075c
0404375c
375c6d72
345c0407
63720273
0276345c
00210f5c
0c8d38c3
c0760296
08040f56
402c1016
303c04eb
094c01c7
8c8c6c00
4ea96c0c
13944007
001c700c
011c7100
4c0b0002
0057123c
0a7c5cbc
0427045c
0404345c
345c6d72
00730407
648d6006
08040856
402c1016
303c04eb
294c01c7
8c8c6c80
6ea96c0c
12946027
001c700c
011c7100
4c0b0002
0057123c
0a7c5cbc
0427045c
0404345c
345c6d72
08560407
00000804
31c3ff96
4c4c240c
042d0809
21c32c89
40374025
00010f5c
01960c8d
00000804
402c1016
303c04eb
294c01c7
8c8c6c80
001c700c
011c7100
4c0b0002
0057123c
0a7c5cbc
0427045c
0404345c
345c6d72
08560407
00000804
402c3016
303c04eb
294c01c7
8c8c6c80
6c0cb0cc
40074ea9
055c1e94
30c30273
fffd341c
0276355c
001c700c
011c7100
4c0b0002
0057123c
0a7c5cbc
0427045c
0404345c
345c6d72
355c0407
63720273
0276355c
345c6006
0c5602bd
00000804
fd967016
402c51c3
14eb292c
01c7303c
6f00c94c
540c8c8c
05897489
033c082d
00b70010
00413f5c
c9c1c74b
0020633c
6f5cc077
076b0021
345c0b41
60270231
60060594
0235345c
700c0253
7100001c
0002011c
123c4c0b
5cbc0057
045c0a7c
345c0427
6d720404
0407345c
0020063c
2f5c0037
548d0001
0e560396
00000804
31c3ff96
4c0c2489
082d0d89
0010013c
2f5c0037
4c8d0001
08040196
00000804
fc967016
402c51c3
303c04eb
294c01c7
8c8c6c80
1489340c
345c504c
68720404
0407345c
315c682b
303c000e
60f70020
00613f5c
c5c1c86b
0020633c
3f5cc0b7
080b0041
033c05c1
00770020
00216f5c
6741684b
001c700c
011c7100
4c0b0002
0057123c
0a7c5cbc
0427045c
0404345c
345c6d72
063c0407
00370020
00011f5c
0496348d
08040e56
fc963016
a48941c3
04eb402c
01c7303c
6c80294c
2c4c6c8c
642b500c
000e325c
0020353c
3f5c60f7
a46b0061
533ca9c1
a0b70020
00413f5c
09c1040b
0020033c
3f5c0077
a44b0021
133ca9c1
20370020
00012f5c
0496508d
08040c56
0136f016
51c3fa96
24eb402c
01c7313c
6f00c94c
8c8c2c0c
540c108c
e0097489
841c87c3
8f5c0007
6f5c00a7
c82d00a1
0010833c
00878f5c
00816f5c
63326009
0074833c
00678f5c
00613f5c
66a96b21
60274089
12c30894
20b72072
00412f5c
00f3408d
617232c3
7f5c6077
e08d0021
001c700c
011c5a00
2c0b0262
0a7c5cbc
0427045c
0404345c
345c6d72
263c0407
40370010
00013f5c
0696748d
0f568076
00000804
f996f016
402c51c3
303c04eb
294c01c7
8c8c6c80
140c308c
41b75489
cea96c0c
3c94c007
323c4489
60070084
43923754
7f5c4177
e48d00a1
32c34409
0007341c
6f5c6137
c02d0081
27c3e197
40f74025
00612f5c
63326409
0074733c
3f5ce0b7
61210041
0010723c
0f5ce077
01b70021
44724489
3f5c4037
648d0001
001c700c
011c5a00
2c0b0262
0a7c5cbc
0427045c
0404345c
345c6d72
6f5c0407
d48d00c1
0f560796
00000804
fc96f016
51c360c3
04eb402c
01c7303c
6c80294c
0c8c2c0c
940c408c
60f77489
602766a9
305c3d94
69720404
0407305c
e006680c
ffff711c
66d23783
cceb7a0c
0393705c
686e7b80
102d0849
63c360d7
c0b7c025
00413f5c
f1a1e869
0010633c
0f5cc077
680c0021
711ce006
3783ffff
660966f2
c629684d
0153c86d
e4f2e849
684d6609
c86900b3
e629c3f2
286be86d
303c3041
60370020
00016f5c
7f5cc0f7
f48d0061
0f560496
00000804
0336f016
50c3fd96
62c371c3
802c6364
25cc50ec
60776409
00213f5c
005d3f5c
935c620c
60570061
98e483c3
323c0635
26c33a1d
01733664
4006706c
00052f5c
20e68cec
3f3c26c3
466400b0
6c6c758c
17c305c3
00063664
c0760396
08040f56
0336f016
01c370c3
636462c3
363cbc2c
354c01c7
15306c80
6c0c2c8c
40074ea9
40c33394
053e243c
0393315c
215423e4
341c69a0
331cffff
1bd47ffe
4029642c
402b4d0d
404b4c6e
406b4c0e
408b4c2e
4c4e4312
315c700b
315c03a6
60720404
0407315c
47cb18c3
602532c3
019367ce
0404315c
315c6572
746c0407
07c36d8c
450616c3
c0763664
08040f56
0136f016
41c370c3
636462c3
363ca02c
154c01c7
4c8c6c00
2ea96c0c
29942007
013c14c3
325c033e
03e40393
61a01654
ffff341c
7ffe331c
345c10d4
6a6f000c
025c10a9
640b0285
0386325c
0404325c
325c6172
02530407
0404325c
325c6572
746c0407
07c36d8c
450616c3
00d33664
0004f524
00040004
80760013
08040f56
236430c3
f5240e24
323c2c2c
454c01c7
6c8c6d00
0444335c
0008341c
f52466f2
00040004
00130004
4004303c
f32462d2
00000804
ff967016
536452c3
353c402c
294c01c7
2c8c6c80
6c0c84cc
60276ea9
60061e94
0427315c
0404315c
315c6d92
c0060407
2006d20f
0225145c
022f645c
145c61c3
2066024d
0276145c
6f5c686c
8cec0005
25c320c6
46646006
0e560196
00000804
fd961016
802c2364
01c7323c
6c80314c
6c0c2c8c
60b76ea9
13946007
135c64cc
21720251
1f5c2077
135c0021
706c0255
00411f5c
00051f5c
21668cec
46646097
08560396
00000804
0136f016
80c3ff96
736472c3
373cc02c
594c01c7
648c2d00
4006accc
02bd235c
235c4006
235c0427
4d920404
0407235c
6ea9640c
1f946027
355c6006
786c0276
2f5c4006
8cec0005
27c32166
46646006
0251255c
341c32c3
60070002
786c1354
2f5c4006
8cec0005
206608c3
600627c3
01134664
0273255c
341c32c3
355cfffe
01960276
0f568076
00000804
fe967016
536452c3
353c402c
894c01c7
8c8c6e00
cdeb6c0c
345c6429
642b0376
0356345c
345c644b
345c0366
61720444
0447345c
145c2006
345c0427
6d920404
0407345c
0464145c
0024313c
31c36cd2
345c6192
684c0467
16c38c8c
600625c3
03334664
0484345c
0024133c
26d22077
6c0c68ac
366415c3
602601d3
0235345c
4f5c686c
4f5c0021
8cec0005
25c32186
46646057
0e560296
00000804
ff963016
802c2364
01c7323c
6e80b14c
6c6c6c8c
000b515c
515cac0e
ac4e001b
002b515c
515cac2e
ac6e003b
2006706c
00051f5c
22a68cec
46646006
0c560196
00000804
0336f016
41c390c3
836482c3
383ce02c
5d4c01c7
cc0c6d00
046c2c8c
215ca44c
323c0404
60071004
60063654
0427315c
deff301c
215c2383
245c0407
400e000b
001b345c
245c604e
402e002b
003b345c
742b606e
04356367
7a4d6026
40060073
215c5a4d
323c0464
66d20404
669232c3
0467315c
215c0153
323c0484
65d20084
639232c3
0487315c
6c4c7c4c
18c309c3
36644006
0f56c076
00000804
0736f016
a0c3fa96
536452c3
1870c02c
01c7353c
6d00594c
ec8c4c0c
64299c8c
702993c3
9f5c93a3
3f5c00a7
702d00a1
933c6449
9f5c1cac
1f5c0087
302d0081
60276aa9
70893e94
941c93c3
19c30001
446628d2
00052f5c
8cec38c3
07b321a6
0404375c
0024733c
2546ead2
00051f5c
88ec28c3
25c321a6
063339c3
4004233c
4ad240f7
3f5c6546
18c30005
21a684ec
37c325c3
78ac0493
15c36c2c
50893664
40b74272
00413f5c
1f5c708d
1f5c0061
28c30005
0ac388ec
25c32306
01f360d7
63727089
1f5c6077
308d0021
2f5c4006
38c30005
22e68cec
600625c3
06964664
0f56e076
00000804
0336f016
80c3fb96
62c371c3
a02c6364
363c3470
554c01c7
2c0c6d00
8c8c6c8c
235c4006
235c0427
4d920404
0407235c
602766a9
50893094
0014323c
2b546007
40f74092
00613f5c
5c29708d
502932c3
613732a3
00813f5c
4117702d
5c4932c3
19ac323c
3f5c60b7
702d0041
6c2c74ac
366416c3
45725089
3f5c4077
708d0021
2f5c4006
39c30005
08c38cec
26c32306
46646006
c0760596
08040f56
ff963016
236441c3
323c202c
454c01c7
0c0c6d00
448c2c8c
600762a9
315c3994
315c0427
6d920404
0407315c
53c36889
00fd541c
3f5ca037
688d0001
a86db029
684d7049
001b545c
680ca86e
411c8006
3483ffff
a20966f2
6229a84d
0153686d
84f28849
a84da209
686900b3
822963f2
315c886d
69720404
0407315c
0484215c
0104323c
32c365d2
315c6492
01960487
08040c56
ff963016
602c51c3
20066c6c
00051f5c
20e68cec
466435c3
0c560196
00000804
31c3ff96
40093264
125440a7
04b440a7
1e944067
40e70093
02331bb4
233c33c4
6046f88c
60376d20
00012f5c
60270093
40860494
0193400d
00f36026
67d22046
60272026
60860494
0053600d
0196200d
00000804
226421c3
31c32009
0004341c
323c6dd2
68070c04
61060494
00d3600d
0080331c
40860394
0804400d
ff96f016
72c360c3
a02c7364
01c7373c
6d00554c
6c0c8c8c
60276ea9
043c1694
20250610
b0bc4106
345c08cb
60720444
0447345c
4006746c
00052f5c
06c38cec
27c32126
46646006
0f560196
00000804
60c3f016
736472c3
373ca02c
554c01c7
8c8c6d00
345c6006
345c0427
6d920404
0407345c
0610043c
41062025
08cbb0bc
0444345c
345c6072
744c0447
06c36c2c
400617c3
245c3664
323c0464
66d20014
609232c3
0467345c
345c0173
341c0484
66d20004
6c0c74ac
17c306c3
0f563664
00000804
fe967016
62c350c3
802c6364
01c7363c
6d00514c
6c0c0c8c
60776ea9
16946007
0484305c
305c6572
0c250487
41062025
08cbb0bc
2f5c706c
2f5c0021
8cec0005
212605c3
605726c3
02964664
08040e56
71c3f016
202c2364
01c7323c
6d00454c
94ccac8c
043cc44c
173c0100
41060010
08cbb0bc
004c375c
d8cc70ef
0300043c
0200143c
0080243c
0180343c
740c6664
7100001c
0002011c
123c4c0b
5cbc0057
055c0a7c
355c0427
6d720404
0407355c
0273345c
345c6272
0f560276
00000804
0336f016
70c3fd96
92c341c3
402c9364
01c7393c
2e80a94c
648cc92c
0870accc
6ea9640c
600760b7
265c4b94
32c30121
0001341c
3c546007
0251355c
60776072
00212f5c
0255255c
000c345c
245c740f
542f002c
004b345c
0266355c
0080053c
00b0143c
b0bc4106
7dac08cb
01066c2c
0100153c
36644046
009c245c
7dac54cf
00866c2c
01c0153c
36644046
00413f5c
00053f5c
88ec28c3
208607c3
609729c3
355c4664
63720273
0276355c
a3460253
00055f5c
88ec28c3
29c321a6
64860133
00053f5c
94ec58c3
29c321a6
46646006
c0760396
08040f56
ff961016
440c41c3
6d2c602c
0010023c
0240133c
b0bc4106
508908cb
610532c3
2f5c6037
508d0001
08560196
00000804
ff963016
402c41c3
10eb292c
01c7303c
6c00094c
100cac8c
6ea96c0c
1f946027
24850025
b0bc4106
708908cb
010503c3
2f5c0037
508d0001
001c740c
011c7100
4c0b0002
0057123c
0a7c5cbc
0427055c
0404355c
355c6d72
00730407
708d6006
0c560196
00000804
0336f016
80c3fe96
72c391c3
c02c7364
01c7373c
ac80394c
30cc948c
0251215c
0014323c
40926ed2
2f5c4077
215c0021
740c0255
39c32deb
60064c29
0946e4bc
0464145c
0804313c
23546007
0889508c
341c30c3
60070002
60061c54
0427345c
0404345c
345c6d92
31c30407
345c6792
88890467
041c04c3
003700fd
00011f5c
784c288d
08c36c6c
49c317c3
36645029
c0760296
08040f56
0136f016
61c3ff96
e92c402c
313c24eb
294c01c7
ac8c6c80
0021865c
433c780c
04c30010
9cbc2106
04c308cb
0240173c
b0bc4106
740c08cb
7100001c
0002011c
123c4c0b
5cbc0057
055c0a7c
355c0427
6d720404
0407355c
0080183c
2f5c2037
588d0001
80760196
08040f56
42c33016
426453c3
301c400b
311c988c
4c0e4103
6045402b
001c4c0e
011c9886
600b4103
07f4213c
ff80341c
400e23a3
10948007
009c301c
4107311c
4000201c
201c4c0e
211c9880
680b4103
fffb341c
618601d3
4107311c
4000201c
201c4c0e
211c9880
680b4103
62723364
540b680e
311c6706
4c0e4107
64c55449
0c564c0e
00000804
40060364
4107211c
341c680b
303c003f
336431ac
301c680e
311c009a
201c4107
4c0ef000
100c303c
f000341c
211c4446
680e4107
00000804
ff961016
618c1364
67c60c8c
2100311c
433c6c0b
60860014
80076037
400f2194
0010313c
7ffe201c
f3ff211c
201c3283
211cc000
32a30c00
20c3604f
301c2364
311c0092
4c0e2100
808c203c
4c0e6045
311c6746
201c2100
4c0e0081
3f5c8037
03c30001
08560196
00000804
211c4006
680b4140
0008341c
680b65f2
63723364
6406680e
2040311c
4c0e4826
00000804
ff963016
12c341c3
440f400c
25c3a089
007f241c
392c533c
0f5ca037
048d0001
215c500c
702c002f
004f315c
0c560196
00000804
311c6486
41262040
600c4c0e
211c4806
680f2040
680f602c
680f604c
680f606c
211c4506
680b2040
0001341c
64867dd2
2040311c
4c0e4226
40066385
4c0f4c0f
4c0f4c0f
211c4506
680b2040
0001341c
08047dd2
40c33016
323c02c3
2580fff0
00d34006
a5a232c4
4025b121
1bf21fe5
08040c56
0736f016
50c3f296
82c371c3
6f3c93c3
06c30330
40a62006
0891bebc
095808bc
0024a01c
2040a11c
2ac36006
4f3c680e
04c30130
420615c3
09585ebc
00305f3c
18c305c3
5ebc4206
04c30958
095834bc
03804f3c
243c4026
06c3f5de
2f3c19c3
60060240
09581abc
70ee6026
2ac36426
500c680e
311c6586
4c0f2040
6085502c
504c4c0f
4c0f6085
6085506c
740c4c0f
211c4806
680f2040
680f742c
680f744c
680f746c
211c4506
680b2040
0001341c
48867dd2
2040211c
7c0f680c
7c2f680c
7c4f680c
7c6f680c
311c6486
40062040
0e964c0e
0f56e076
00000804
201c0364
211c9880
680b4103
61723364
680b680e
fff7341c
0cf2680e
009c301c
4107311c
4000101c
680b2c0e
fffb341c
61860153
4107311c
4000101c
680b2c0e
62723364
0804680e
326432c3
301c6df2
311c00a0
5fe64107
40ab4c0e
009e301c
4107311c
60270553
301c0d94
311c00a4
5fe64107
40ab4c0e
00a2301c
4107311c
60470393
301c0d94
311c00a8
5fe64107
40ab4c0e
00a6301c
4107311c
606701d3
301c0d94
311c00be
5fe64107
40ab4c0e
00bc301c
4107311c
63464c0e
4107311c
4c0e5fe6
6045408b
21c34c0e
301c2364
311c9888
4c0e4103
808c213c
4c0e6045
6006402b
4107311c
321c4c0e
5fe6009c
404b4c0e
311c6186
4c0e4107
008e321c
4c0e5fe6
6446406b
4107311c
40094c0e
4c0e6785
00000804
22640364
141c2312
65c6fff8
4107311c
33646c0b
0300141d
0044323c
303c66d2
213c1900
0213180c
0084323c
303c66d2
213c17e0
0113080c
0024323c
0280203c
313c65d2
6980088c
68800053
036403c3
00000804
326430c3
05946027
311c6446
00d34107
301c68f2
311c009a
201c4107
4c0e0403
00000804
f996f016
12c331c3
60b73264
0020723c
311c6486
201c2040
4c0e0081
01c04f3c
343c6926
400cf87e
000f245c
4806700c
2040211c
602c680f
002f345c
01c06f3c
fa4e363c
604c680f
004f345c
01c05f3c
fc4e353c
6189680f
00cd3f5c
3f5c6006
3f5c00d5
3f5c0041
0f3c00dd
303c01c0
680ffe4e
0100201c
6409500e
141c13c3
207700e3
00212f5c
00752f5c
345c6006
345c001f
345c003f
4006005f
00dd2f5c
211c4506
680b2040
0001341c
700c7dd2
211c4806
680f2040
680f780c
680f740c
680f600c
85062006
2040411c
027302c3
341c700b
7dd20001
600f7c81
682c5c80
684c600f
686c600f
213c600f
40370100
00011f5c
23c36097
ebb421e4
211c4506
680b2040
0001341c
65867dd2
2040311c
03c36c0c
0f560796
00000804
000620c3
28060a0f
a040111c
323c29cf
698f0340
323c294f
690f0240
0b8f28cf
32c32085
327e133c
32c36b0f
2a7e133c
2a2f6a8f
00000804
fd967016
426442c3
201c600f
211c8010
404f0008
600620c3
633c0353
c0770010
00213f5c
60674205
f5240694
00040004
00130004
601c280f
611c8010
c84f0008
643c2205
c037ff00
00014f5c
e6948007
41806412
351c684c
684f6000
311c69c6
6c0b2100
0001341c
40b74086
13946007
236420c3
0098301c
2100311c
203c4c0e
6045808c
69464c0e
2100311c
0081501c
80b7ac0e
00416f5c
039606c3
08040e56
fd967016
426442c3
201c602f
211c8010
404f0008
600620c3
633c0353
c0770010
00213f5c
60674205
f5240694
00040004
00130004
601c282f
611c8010
c84f0008
643c2205
c037ff00
00014f5c
e6948007
41806412
351c684c
684f6000
311c6bc6
6c0b2100
0001341c
40b74086
13946007
236420c3
009e301c
2100311c
203c4c0e
6045808c
6b464c0e
2100311c
0085501c
80b7ac0e
00416f5c
039606c3
08040e56
fe967016
61c343c3
22646364
602c4037
6586ad2c
4107311c
4c0e4046
73ae60a6
0203245c
311c6486
4c0e4107
301c53eb
311c80b2
4c0e4103
86a4201c
4103211c
3364680b
680e6372
60277269
65c61194
4107311c
13642c0b
6c0b6705
412c3364
203c08c9
69801b0c
0af413e4
3f5c0453
03c30001
094a84bc
00870364
72691a35
07946027
311c6446
201c4107
4c0e0100
311c6446
00264107
321c0c0e
cc0e015e
641276ac
000f351c
400676af
00734077
60776066
00212f5c
029602c3
08040e56
0336f016
50c3fe96
32c381c3
60373264
2130002c
e14c81ac
33abd38b
245c4026
65860165
4107311c
245c2c0e
64860203
4107311c
53eb4c0e
80b2301c
4103311c
201c4c0e
211c86a4
680b4103
63723364
75ec680e
341c6c4c
60070002
618c1754
03a1335c
129460a7
01c7363c
6c8c7d80
235c6ccc
32c30273
0001341c
20c767d2
313c0535
13c3ffc0
383c1364
6ef20014
d2bc28c3
30c30957
68d23264
06946087
0004f524
00040004
72690013
16946027
311c65c6
2c0b4107
67051364
33646c0b
08c9552c
1b0c203c
13e46980
644642d4
4107311c
0101001c
145c05d3
20070149
2f5c2c94
02c30001
094a84bc
00870364
752c3035
001c6c0c
011cff00
308300ff
0100101c
0001111c
32e421c3
74ec1094
0451335c
0b946027
311c6446
20864107
63462c0e
4107311c
4c0e5fe6
311c6446
00264107
00930c0e
145c2006
29c3014d
64126aac
000f351c
60066aaf
00736077
00770066
00211f5c
029601c3
0f56c076
00000804
fe967016
840c448c
680c212c
525c0c0b
a07702f1
0754a027
60076057
60671454
01b33094
303c0c6b
7f32fff0
0020633c
1f5cc037
125c0001
047302f5
325c6086
03f302f5
00215f5c
02f5525c
0404325c
325c6092
c7cb0407
7fe536c3
67ce3164
06156007
0004f524
00040004
60260013
3523b20b
615c33e3
36830253
0256315c
0e560296
00000804
fe967016
212c20c3
838b01ac
01c7343c
6f00c94c
ac8c8c0c
36c3c026
3623d20b
0253615c
315c36a3
60260256
686c622d
655c100c
c5f202d1
153c6dec
00930470
153c6dec
366404c0
255c700c
4c2d0299
c006700c
7389cc0d
10946027
300c514c
808c323c
66ee3203
635c700c
c0720169
2f5cc077
235c0021
92a9016d
85f28037
00013f5c
02c5355c
455c8006
c0060396
02b5655c
02ad655c
0305655c
0e560296
00000804
30c37016
21ac812c
203c078b
cd4c01c7
ac8c6b00
4c0c14cc
ca0b6026
33e33623
0253245c
345c3283
60060256
013d315c
66ed668d
672d670d
c20fc006
0225305c
022f605c
024d305c
02bd355c
08040e56
30c31016
01ac212c
243c838b
8d4c01c7
4c0c6a00
627267eb
301c67ee
311cbed6
694f8e89
5555401c
6aa6884e
800668cd
0856822d
00000804
bed6201c
8e89211c
201c414f
404e5555
40cd4aa6
00000804
20c33016
026401c3
89ac292c
353cb38b
a94c01c7
4c0c6e80
04940047
647267eb
002700b3
67eb0494
67ee6372
dabc02c3
6006095c
0c56722d
00000804
402c1016
878b29ac
02c7343c
4e008a6c
34c388eb
68ee6025
6c29612c
05946027
4f0c60ec
4f0f4025
627266ac
085666af
00000804
72c3f016
400c1364
8cac608c
ac0b6c0c
60a76929
6aa92a94
27946007
353cd02c
62520057
0377333c
128d033c
5cbc2c86
102f0a7c
012c301c
012b031c
201c0b35
353c1388
6352228d
ff6a321c
03e46132
702f0235
70e4102c
f5240634
00040004
00130004
00530320
0f560006
00000804
50c37016
31cc802c
0b8b51ac
02c7303c
0f00d26c
341c6aac
6ad20020
32c344ab
64ae6025
36c3c12b
612e6025
44cb0133
602532c3
c14b64ce
602536c3
708c614e
05c36c2c
36642026
6c6c708c
366405c3
08040e56
ff967016
51c340c3
2f5c4006
60c9001d
21546087
08b46087
11546047
13b46047
2d946027
60c70453
60c70654
60e71a14
03f32694
00402f3c
02137e06
00402f3c
0353caa6
2f5c5e06
201c001d
211ca184
03330013
00402f3c
323c7fe6
0273ffde
00402f3c
0113c006
00402f3c
fed361e6
00402f3c
623cd546
00b3ffde
a084201c
0013211c
204610a9
75ac0233
cca1c809
36c3d0c9
7f327fe5
313c4980
13c30010
303c1364
03c3fff0
00070364
b00fef94
0e560196
00000804
ff963016
602c40c3
618cadcc
1fc36c0c
20173664
30c314a9
668e6045
6c6b70cc
6d004017
6017644f
0100233c
0c6b70cc
65af6800
4c0d54c9
14a965ac
54a90c2d
624532c3
05c3644e
095d80bc
0c560196
00000804
40c31016
41ec61ac
21466c0c
36644849
0948bebc
6c8c702c
04c36c6c
08563664
00000804
0136f016
50c3ff96
9dcce02c
0130ddac
08c340ec
101c600c
111cff00
318300ff
0100001c
0001011c
31e410c3
325c0794
70cd0469
0421025c
202610ad
012d165c
65f2700c
6dcc7c6c
366405c3
680c28c3
ff00001c
00ff011c
500c3083
0100101c
0001111c
30e401c3
29ac0794
400638ef
012d265c
7c8c0353
10a929ac
404520c3
0f5c0046
8c0c0005
600605c3
75ac4664
6c0c55ec
210605c3
36644849
0948bebc
6c6c7c8c
366405c3
80760196
08040f56
0736f016
a1c360c3
e02ca264
bdac1dd0
8e2421f0
0046f524
095edcbc
4004343c
f32462d2
0129355c
04946027
0129355c
355c7ef2
60270131
355c0494
7ef20131
0948b6bc
0001a31c
001c0c94
29c30270
cebc2849
7c8c094b
06c36c4c
02933664
2c0c38c3
798c28d2
06c36c4c
60063664
680f28c3
04e1001c
284929c3
094bcebc
38c34026
e0764d0d
08040f56
410c30c3
6dec080c
66f26c49
311c6306
22064107
602702f3
63060694
4107311c
02132406
07946047
311c6306
101c4107
01130200
07946067
00e0301c
4107311c
2c0e2026
3664682c
00000804
326430c3
634666f2
4107311c
02f34206
06946027
311c6346
44064107
60470213
63460794
4107311c
0200201c
60670113
301c0794
311c00e2
40264107
08044c0e
326430c3
638666f2
4107311c
02f34206
06946027
311c6386
44064107
60470213
63860794
4107311c
0200201c
60670113
301c0794
311c00e4
40264107
08044c0e
226420c3
013e301c
4107311c
00ff101c
301c2c0e
311c013c
4c0e4107
20266105
301c2c0e
311c0142
20064107
61452c0e
61852c0e
0082101c
47f22c0e
311c6306
42064107
03134c0e
06944027
311c6306
24064107
40470213
63060794
4107311c
0200101c
40670113
301c0794
311c00e0
20264107
08042c0e
ff96f016
ccc9612c
08b7463c
3fff441c
2c4961ec
ac4b2037
6c0c61ac
7f5c2006
27c30001
201c3664
211c9880
680b4103
61723364
2017680e
6c062ef2
4107311c
04e1201c
6b064c0e
4107311c
0ce1701c
0633ec0e
21c32017
0b944027
311c6c46
701c4107
ec0e04e1
311c6b46
04134107
32c34017
0d946047
008a301c
4107311c
04e1701c
301cec0e
311c0088
02134107
32c34017
0f946067
00c4301c
4107311c
04e1701c
301cec0e
311c00c2
101c4107
2c0e0ce1
311c6146
40064107
62454c0e
e1cf701c
2017ec0e
406721c3
321c0594
e02600c8
201cec0e
211c9880
680b4103
fff7341c
201c680e
211c0200
680b4107
fffd341c
263c680e
6cc608f7
4107311c
61864c0e
4107311c
2000101c
a0672c0e
321c0854
e8060090
101cec0e
2c0e0200
009c301c
4107311c
0400201c
701c4c0e
ec0e8000
0654a067
40866085
60854c0e
301c4c0e
311c00a8
e0864107
62c5ec0e
6346ec0e
4107311c
0230101c
321c2c0e
402600c8
64464c0e
4107311c
ec0ee806
21c32017
311c6006
e4864107
09544047
21c32017
07944027
311c6006
e2464107
0253ec0e
27f22017
311c6006
40264107
01534c0e
73c36017
0694e067
311c6006
27064107
a0672c0e
60173b54
301c69f2
311c00a4
e0264107
6085ec0e
20170193
402721c3
301c0b94
311c00a0
71c34107
61052c0e
62c5ec0e
20170453
404721c3
301c0e94
311c00a4
e0264107
301cec0e
311c00a0
ec0e4107
023363c5
21c32017
0e944067
00a4301c
4107311c
ec0ee026
00a0301c
4107311c
6105ec0e
61c6ec0e
4107311c
017c101c
40062c0e
4107211c
341c680b
343c003f
336431ac
301c680e
311c009a
201c4107
4c0ef000
3c00441c
100c243c
311c6446
4c0e4107
ea066745
0196ec0e
08040f56
036421c3
301c2264
311c013e
101c4107
2c0e00ff
013c301c
4107311c
20c34c0e
61454b72
08044c0e
036421c3
301c2264
311c013e
101c4107
2c0e00ff
013c301c
4107311c
62054c0e
08040c0e
226421c3
2c0c620c
009e301c
4107311c
15544007
06944027
00a2301c
4107311c
404701d3
301c0694
311c00a6
00f34107
07944067
00bc301c
4107311c
64ae6c0b
311c6386
6c0b4107
6006648e
4107311c
642e6c0b
311c6186
6c0b4107
6bc6644e
4107311c
640d6c0b
311c6446
6c0b4107
0804646e
780c313c
213c2089
001c00f4
011c8000
3083007f
59ac323c
236423c3
190b113c
011a301c
4107311c
301c4c0e
311c0086
2c0e4107
00000804
02c330c3
12643264
29546007
13942027
00ba201c
4107211c
3364680b
680e6772
9880201c
4103211c
101c680b
31a38000
02133364
00ba201c
4107211c
3364680b
680e6e72
98a0201c
4103211c
3364680b
680e6272
0104301c
04b3600e
11942027
00ba201c
4107211c
341c680b
680eff7f
9880201c
4103211c
341c680b
02137fff
00ba201c
4107211c
341c680b
680ebfff
98a0201c
4103211c
341c680b
680efffb
200e2546
00000804
30c31016
13643264
180c013c
0e546047
04b46047
18946027
608700d3
61070b54
01b31394
0280303c
303c0293
6505088c
313c0213
321c300c
01730190
200c313c
017e321c
f52400d3
00040004
00130004
0856680e
00000804
41c31016
213c200c
301c808c
311c98ae
4c0e4103
236421c3
4c0e6045
213c202c
301c808c
311c9888
4c0e4103
236421c3
4c0e6045
213c204c
6245808c
21c34c0e
60452364
206c4c0e
808c213c
9898301c
4103311c
21c34c0e
60452364
500b4c0e
4c0e66c5
6045502b
08564c0e
00000804
42c31016
323c4009
60070024
201c1154
211c9884
680b4103
fff7341c
680b680e
fffb341c
680b680e
61723364
323c07f3
60070044
201c1154
211c9884
680b4103
fffd341c
680b680e
fff7341c
680b680e
62723364
323c0293
60070084
201c1654
211c9884
680b4103
fffd341c
680b680e
fffb341c
680b680e
63723364
01c3680e
90bc14c3
02730961
600d6026
9884201c
4103211c
341c680b
680efffd
341c680b
680efff7
341c680b
680efffb
08040856
988c301c
4103311c
33646c0b
988e201c
4103211c
113c280b
301c81ac
311c98b6
4c0b4103
60452364
333c6c0b
0006812c
e0bf201c
12833283
025431e4
08040026
1364ff96
0161205c
301c4512
311c02aa
4c0e4107
6085402b
404b4c0e
4c0e6045
6b1260c9
236423c3
02ac301c
4107311c
67054c0e
42eb2c0e
4c0e6045
0169105c
0024313c
301c69d2
311c02e8
4c0b4107
41722364
313c4c0e
69d20044
02e8301c
4107311c
23644c0b
4c0e4272
02e8301c
4107311c
23644c0b
4c0e4072
680b23c3
4000341c
301c7dd2
311c02e8
0c0b4107
320b303c
2f5c6037
02c30001
08040196
42c33016
526450c3
33641364
013e201c
4107211c
00ff001c
201c080e
211c013c
a80e4107
036404c3
080e4105
808c043c
0142201c
4107211c
4145080e
301c680e
311c0158
201c4107
4c0e0082
0140301c
4107311c
63062c0e
4107311c
a0070206
63061554
4107311c
a0270406
63060f54
4107311c
0200001c
0854a047
0794a067
00e0301c
4107311c
0c0e0026
08040c56
fe967016
41c352c3
67c64364
2100311c
341c6c0b
13c30001
40774086
1d546007
313c0753
4180200c
180c313c
cc0c7580
cc4bc80f
602536c3
3ffe601c
0001611c
601c3683
611c8000
36a30c00
313c684f
60370010
00011f5c
336431c3
e21434e4
200c313c
41807e05
6e72684c
20c3684f
301c2364
311c0092
4c0e2100
808c203c
4c0e6045
311c6746
201c2100
4c0e0081
60776006
00216f5c
029606c3
08040e56
ff963016
526451c3
40372264
8ccc608c
094c56bc
0200043c
094c78bc
010c201c
4107211c
3364680b
680e6072
0694a027
133c34c3
4145204e
aff20133
133c34c3
201c22ce
211c0116
280f4107
3f5c03c3
13c30001
0960f4bc
301c50cc
311c010e
4c0f4107
608550ec
01964c0f
08040c56
ff963016
602c50c3
01f38d2c
6265558c
480c6212
318005c3
51c92664
602532c3
2f5c6037
51cd0001
602771c9
0196f035
08040c56
63ae6006
080463ee
41c31016
22644364
2d2c602c
18544007
0ce9620c
336430c3
0c9443e4
30236026
215c33e3
32830243
0236315c
315c6006
60260246
215c3423
32a30243
602600f3
33e33423
0243215c
315c3283
08560246
00000804
0736f016
51c3a0c3
936492c3
28c30030
840cc9ac
66f239c3
0004f524
00040004
648c0013
02f1335c
6047e006
05b32694
335c748c
602702f1
f5240694
00040004
00130004
60a77129
28c30794
6dac686c
320b0ac3
73893664
6027100c
748c0794
0393135c
096240bc
86bc0073
1a4d0967
0010373c
736473c3
db1479e4
510d5a49
58bc1a49
10ed0967
4026748c
02c5235c
0f56e076
00000804
31c33016
8c8c240c
0383245c
0393545c
602535c3
189423e4
4f8b61ac
02c7323c
4e80a26c
30c30a6b
6a6e6025
143c040c
10bc04c0
40260967
02d5245c
0404345c
345c6192
0c560407
00000804
e6bc2126
08040949
f8bc2126
08040949
0336f016
80c3f896
e02c61c3
648c9d2c
2410ac0c
00400f3c
43862006
0891bebc
325c588c
60720404
0407325c
31c333cb
73ce6025
32c353eb
0002341c
7d4c6ad2
6c0c6c8c
3f5c6c0b
3f5c0096
00f300a6
3f5c740b
340b0096
00a61f5c
2f5c542b
744b00b6
3f5c6332
7c6c00c6
08c38d6c
2f3c2046
36c30040
7c6c4664
460b19c3
1f5c2006
8cec0005
600608c3
08964664
0f56c076
00000804
6d2c602c
08040feb
40c31016
f8bc24ab
702c0949
40066d2c
08564e0d
00000804
40c31016
e6bc24ab
702c0949
40266d2c
08564e0d
00000804
41c31016
096472bc
98bc04c3
085608c9
00000804
0736f016
91c380c3
8ebc52c3
70c30895
64c39fe6
0001a01c
05c30333
08ce0cbc
28c30364
333c680c
6fa00e1d
05156007
616460c3
01938086
043543e4
616460c3
3a3c43c3
33e3000d
a0075383
39c3e794
06c38c0f
0f56e076
00000804
8e241016
402cf524
096494bc
343c0164
62d24004
0856f324
00000804
ff961016
7fe640c3
602c6037
00ab6ad2
089580bc
05f20037
1fc304c3
0964c2bc
01960017
08040856
fc967016
61c340c3
40772264
536453c3
4d2c602c
600769c9
133c1154
2037fff0
00013f5c
0f5c60b7
09cd0041
31c32097
023c6265
00f73a1d
618c00d3
1f3c6c0c
366400c0
202660d7
6c4f2f2e
235c4006
af4e01e5
086950cc
420520c3
1f5c4d00
123c0021
780f00df
049602c3
08040e56
fe967016
61c350c3
40372264
436443c3
6c0c618c
00401f3c
60573664
2f2e2026
40066c4f
01e5235c
54cc8f4e
21c32869
4d004205
00011f5c
00df123c
02c3780f
0e560296
00000804
226420c3
323c1364
64d20014
180c313c
323c02b3
64d20044
300c313c
323c00d3
66d20084
200c313c
0240321c
323c0133
03c30024
313c67d2
321c100c
03c300c8
08040364
13647016
313c402c
294c01c7
708c8c80
cc6cac4c
2f0b692c
133c35c3
500c026f
21250a09
64bc23c3
301c0961
742e00fb
0e29700c
0104101c
0060253c
096164bc
580e4366
0148301c
582e784e
0e56786e
00000804
fd963016
644c51c3
0100233c
2c6960cc
602c8880
50092d2c
241c4077
4037000f
00013f5c
29b460c7
233c6026
323c200d
60070554
323c1494
60070024
3f5c1e54
30640021
0060013c
02156007
143c01c3
88bc0080
30c30942
6ff23264
355c6006
100901e5
2026102d
d6bc300d
045c0949
4006013f
007340b7
60b76026
00411f5c
039601c3
08040c56
0336f016
70c3f996
c02c81c3
99acb92c
303c138b
594c01c7
6c4c6d00
60262c69
012d345c
0131345c
300c313c
0035233c
2f5c40b7
20640041
0c0938c3
941c90c3
393c0040
6077092c
00210f5c
00750f5c
2f5c4186
0f3c007d
20270100
15c30394
153c0073
82bc0060
5f3c0942
0f3c00e0
183c0160
82bc0020
b0ef0942
0c497dec
095edcbc
0006788c
00050f5c
07c38c0c
41c615c3
46646026
c0760796
08040f56
0f36f016
a0c3fc96
3db0e02c
478b19c3
313c12c3
5d4c01c7
7810cd00
788cb86c
20260c10
135c39c3
335c012d
618c0131
1f3c6c0c
366400c0
423c40d7
74890020
14496712
31ac103c
0055013c
3f5c00b7
680d0041
082d0446
035c7d2c
30c30129
0040341c
013c67d2
00770255
00211f5c
5449280d
7d2c46f2
133c04c3
00b30060
04c3788c
0400133c
b0bc40c6
043c08cb
1b3c0060
40c60160
08cbb0bc
4f8b39c3
033c7dec
106f2a1d
0100043c
00401b3c
b0bc4066
18c308cb
326d2509
6c0c7c6c
16c30ac3
03643664
086e28c3
f52406f2
00040004
00130004
38c3114e
716e6c0b
002b08c3
18c3118e
6332644b
388c71ae
01c0043c
02d1215c
28e543f2
29850053
b0bc40a6
788c08cb
0299035c
010d045c
65ec1ac3
dcbc0c49
60d7095e
68ef29c3
00067c8c
00050f5c
0ac38c0c
448620d7
46646026
f0760496
08040f56
fb96f016
802c70c3
b1ac512c
2d09620c
01c7313c
6c80314c
603c0c2c
602604f0
012d355c
0131355c
12c36149
20c562f2
62726612
2f5c60f7
205c0061
305c027d
23c30271
40b740c5
00413f5c
2f5c6137
205c0081
063c0285
40c60020
08cbb0bc
708cd4ef
21c32117
40774045
00212f5c
1f5c2006
8c0c0005
16c307c3
46646026
0f560596
00000804
40c31016
12c301c3
36bc48d2
712c0943
2d090066
0872a2bc
08040856
fb961016
323c21c3
43c3021e
001f441c
3f5c8077
680d0021
405c840c
68090017
640c60cd
06947fe7
63e76809
64a60394
80060573
813780f7
00812f5c
433240b7
34c38117
0007341c
343c8522
341c308d
6bd20001
610040d7
00414f5c
40258ced
4f5c4037
80f70001
32c34117
61376025
e39464a7
46f240d7
0004f524
00040004
3f5c0013
305c0061
05960165
08040856
20c3fc96
44a72264
61862354
44c760f7
40f72154
1e5444e7
07b44147
0010123c
3f5c20b7
01b30041
ff50323c
3f5c6077
63270021
123c08b4
20370020
00013f5c
011360f7
0004f524
00040004
20060013
3f5c20f7
03c30061
08040496
fe961016
200940c3
05004029
6ebc24a6
00370a7c
00013f5c
1f5c6077
300d0021
51806332
31c32057
0007341c
313c2849
341c308d
6af20001
12c34057
0161245c
3120341d
6ce97180
3f5c6077
03c30021
08560296
00000804
ff961016
326430c3
22641264
088c433c
40278037
40472254
27f21894
0001361c
0014133c
03332037
0a942027
0006341c
0002361c
7f327fe5
603769a0
f52401d3
00040004
00130004
40672037
f5240654
00040004
00130004
00011f5c
019601c3
08040856
fc961016
423c2264
8077ffc0
00213f5c
38356027
24944047
688b402c
17946027
03b9325c
13946027
0259325c
8a4960b7
03c3025c
6ebc13c3
00370a7c
4f5c04c3
14c30001
00413f5c
00d323c3
125c0a49
225c03b1
b2bc0259
02640967
40270113
604c0494
00730ca9
0c29606c
20f724a6
303c0fd2
7fe50016
f88c233c
6d2064e6
01c300d3
096786bc
326430c3
3f5c60f7
03c30061
08560496
00000804
30c3ff96
333c3264
7932080d
60376072
00013f5c
019603c3
00000804
0f36f016
60c3ff96
a3c382c3
726471c3
19c32030
4006a52c
6e244037
f524b3c3
648c1ac3
8c0ce3f2
8c2c0053
43d257ab
1754e007
6c2c79ac
1fc30046
366420c3
650b18c3
32e444eb
6d200754
00031f5c
3130341d
700e6980
255c500b
00930226
0223355c
7a0c700e
310d2d69
0954e027
646c19c3
06c36c0c
36641ac3
0073106e
506e500b
654b18c3
704e6312
502e452b
40043b3c
f32462d2
f0760196
08040f56
0736f016
30c3fd96
003091c3
0020513c
21ac08c3
6ce96e0c
333c678e
414c01c7
980ccd00
ec0c788c
72ad6006
120e078b
39c3586c
a0c30c09
0040a41c
310c3a3c
0f5c60b7
088d0041
526d4026
201c678b
63d20108
487223c3
043c51ee
15c30160
094282bc
7c0e756b
1c2e158b
631275ab
18c37c4e
235c652c
32c30129
0040341c
09c369d2
31c32009
0020341c
402663d2
746c538d
150b714f
3649104e
566930cd
754b5d0d
788c7c6e
035c0026
788c02d5
04c0033c
01c0153c
b0bc40a6
788c08cb
0109155c
241c21c3
4077001f
00210f5c
029d035c
555c788c
a5320109
1f5ca037
135c0001
0396028d
0f56e076
00000804
0336f016
40c3f596
52c391c3
01408f3c
200608c3
bebc4206
7f3c0891
07c30040
42062006
0891bebc
42774006
702c42b7
39c3cc4c
a6f262d2
0004f524
00040004
71ac0013
00666c2c
404618c3
2f5c3664
32c300b1
003f341c
60376672
00013f5c
00b53f5c
09c398cc
28c317c3
02403f3c
78ec4664
220607c3
2f5c3664
540d0021
00293f5c
2f5c742d
544d0031
00a13f5c
2f5c746d
548d00a9
00b13f5c
000674ad
c0760b96
08040f56
4d49620c
0006440d
00000804
fe961016
23c36009
10546007
284c402c
133c202f
2037fff0
00013f5c
4f5c6077
800d0021
604f63f2
02c3602f
08560296
00000804
4006ff96
6009444f
204f64f2
0093202f
2c4f604c
4009204f
602532c3
2f5c6037
400d0001
08040196
ff963016
602c52c3
620c8d6c
6d495309
103423e4
631272e9
0d00504c
40c615c3
08cbb0bc
13c37309
20372025
00012f5c
0196530d
08040c56
ff961016
602c10c3
12e98d6c
6d49660c
103530e4
180c303c
0c80302c
40c612c3
08cbb0bc
32c352e9
60376025
00011f5c
019632ed
08040856
fe967016
a16c62c3
02338006
180c343c
0d00544c
40c616c3
08cbeabc
007703f2
243c0193
40370010
00014f5c
34e47709
201ceeb4
407700ff
00213f5c
029603c3
08040e56
fe967016
a16c62c3
02338006
180c343c
0d00542c
40c616c3
08cbeabc
007703f2
243c0193
40370010
00014f5c
34e476e9
201ceeb4
407700ff
00213f5c
029603c3
08040e56
f896f016
61c340c3
726472c3
01000f3c
42062006
0891bebc
ad6c702c
5689720c
20066d49
41c320f7
4a1423e4
740c0a53
243c6e00
2c090280
3a942007
4c0d4026
6e00740c
123c26c3
2c2d009f
6e00740c
0020033c
40c612c3
08cbb0bc
6e00740c
0080033c
0070163c
b0bc4206
740c08cb
033c6e00
163c0180
42060170
08cbb0bc
6e00740c
0180033c
01001f3c
eabc4206
04d208cb
00612f5c
768956ad
202513c3
2f5c2077
568d0021
60b76006
20d70293
602531c3
1f5c6037
20f70001
40d742c3
37e432c3
f524b514
00040004
00130004
20b720e6
00412f5c
089602c3
08040f56
fa967016
61c340c3
5f3c6264
05c30080
42062006
0891bebc
40774006
70090293
09946027
0180043c
420615c3
08cbeabc
10940007
23c36057
40374025
00013f5c
85056077
32c34057
ea1436e4
00ff301c
2f5c6077
02c30021
0e560696
00000804
0736f016
50c3f396
126442c3
9f3c2037
09c30190
42062006
0891bebc
0310af3c
20060ac3
bebc4066
6f3c0891
06c30090
42062006
0891bebc
02908f3c
200608c3
bebc4106
742c0891
ec4cad6c
1f5c3009
5029018d
01952f5c
3f5c7049
3069019d
00cd1f5c
2f5c5089
70a900d5
00dd3f5c
2f5c140c
12c30001
096a7cbc
326430c3
21c32017
193432e4
0287333c
0c80340c
60276009
9ccc1294
16c30305
38c329c3
7cec4664
220606c3
0ac33664
406616c3
08cbeabc
04d20077
00ff101c
2f5c2077
02c30021
e0760d96
08040f56
1f36f016
90c3f396
43c3a1c3
c264c2c3
01908f3c
200608c3
bebc4206
bf3c0891
0bc30310
40662006
0891bebc
00906f3c
200606c3
bebc4206
5f3c0891
05c30290
41062006
0891bebc
682c29c3
70092c50
018d3f5c
2f5c5029
70490195
019d3f5c
2f5c5069
708900cd
00d53f5c
2f5c50a9
7ac300dd
60776006
0413abc3
60277c09
39c31594
073c8ccc
16c30080
35c328c3
29c34664
06c368ec
36642206
16c30ac3
eabc4066
000708cb
60571054
402523c3
3f5c4037
60770001
4057e505
3ce432c3
301cde14
607700ff
00212f5c
0d9602c3
0f56f876
00000804
602c1016
620c8d6c
4d49100c
0287123c
08cb9cbc
728d6006
085603c3
00000804
30c3f016
808c603c
40c30006
53c310c3
e1e65364
110d353c
341c5ca0
32230001
03c330a3
363c0364
341c110d
32230001
43c334a3
20254364
ed942207
802c043c
08040f56
0336f016
90c3fc96
800651c3
807774c3
80f784c3
40d7c3c6
208d393c
0f5c6037
3f5c0001
61e70061
605714b4
270323c3
3f5c4077
13c30021
34031003
230320c3
0001241c
0014313c
09ac323c
83a33623
23c360d7
40f74025
4407dfc5
e0770654
403c74c3
fb130014
e0b7e006
653c3c06
453c00c0
053c0080
40970040
208d383c
0001341c
62f24186
3f5c4066
60e70041
609709b4
323c6212
540c300d
740f32a3
61e70353
323c07b4
400c100d
600f32a3
62e70253
313c09b4
323cfe00
500c300d
700f32a3
313c0113
323cfc00
f80c300d
780f37a3
32c34097
60b76025
64072085
140ccd94
096b8ebc
45c3140f
024e043c
096b8ebc
45c3100f
044e043c
096b8ebc
45c3100f
064e043c
096b8ebc
0496100f
0f56c076
00000804
fe963016
436441c3
620c202c
40060c29
a0574077
01c7353c
6d00454c
69eb4c0c
0a9434e4
60276a89
6a690794
04946027
00213f5c
a0570173
602535c3
60773364
e83530e4
00ff501c
603735c3
00012f5c
029602c3
08040c56
c0963016
4d2c602c
10003f3c
533ca006
ab8b805e
000e535c
0161525c
001d5f5c
886c414c
60862fc3
40964664
08040c56
c0963016
620c802c
353cad09
b14c01c7
6c2c6e80
4f5c8006
ae890005
000d5f5c
8c6c614c
60462fc3
40964664
08040c56
c0967016
61c340c3
602c6364
6c2c6c6c
36642869
10002f3c
805e023c
ac6c714c
16c304c3
60262fc3
40965664
08040e56
bf967016
61c350c3
202c6364
8feb652c
341c34c3
81860024
69f28037
6c4c646c
48892869
30c33664
60373264
10403f3c
00012f5c
805e233c
886c554c
16c305c3
602623c3
41964664
08040e56
bf967016
61c350c3
402c6364
6da9692c
20372186
07946027
6c8c686c
30c33664
60373264
10403f3c
00012f5c
805e233c
886c554c
16c305c3
602623c3
60174664
742c6af2
6d8c4c4c
05c3880c
03b3135c
46644046
0e564196
00000804
c0961016
3f5c6006
620c0005
4f5c8d29
614c000d
2fc38c6c
46646046
08564096
00000804
b896f016
42c360c3
736471c3
744ca02c
125c6d8c
3664001b
126410c3
00ff131c
313c2a54
554c01c7
6c0c6d00
002b245c
08962f5c
003b245c
08a62f5c
004b245c
08b62f5c
005b245c
08c62f5c
006b245c
08d62f5c
007b245c
08e62f5c
60276ea9
746c0a94
06c36ccc
10402f3c
30c33664
00533264
60376186
00012f5c
00252f5c
8c8c794c
17c306c3
00402f3c
46646026
0f564896
00000804
0136f016
70c3bf96
836481c3
952ca02c
6d8c744c
001b125c
60c33664
40466264
631c4037
135400ff
01c7363c
6d00554c
6ea96c0c
09546027
0121245c
341c32c3
82260008
63d28037
40374006
10403f3c
00014f5c
805e433c
888c5d4c
18c307c3
602623c3
40174664
18944007
01c7363c
6e00954c
335c6c8c
341c0444
544c0001
682c69d2
16c307c3
00014f5c
366424c3
68ac00b3
16c307c3
41963664
0f568076
00000804
0136f016
60c3b296
81c342c3
e02c8364
10005f3c
200605c3
bebc4206
20060891
33773337
13802f3c
001c345c
f47e323c
003c145c
345c282f
684f005c
007c145c
3f3c286f
145c1380
133c009c
145cec7e
2c2f00bc
00dc145c
145c2c4f
2c6f00fc
84cc3c4c
15c302c3
3f3c23c3
46641300
6cec7c4c
220605c3
60063664
00053f5c
340c2fc3
000f125c
325c742c
344c002f
004f125c
325c746c
794c006f
06c38c6c
622618c3
4e964664
0f568076
00000804
bf96f016
42c360c3
736471c3
744ca02c
125c6d8c
3664001b
126410c3
00370046
00ff131c
313c2954
154c01c7
680c4c00
01866ea9
60270037
688c1f94
245c6ccc
4c0f002c
004c045c
245c0c2f
235c006b
045c0266
0d8f007c
009c245c
045c4daf
0dcf00bc
00dc245c
744c4def
06c36d0c
60063664
3f3c6037
0f5c1040
033c0001
594c805e
06c3888c
23c317c3
46646026
0f564196
00000804
0336f016
60c3bf96
81c342c3
a02c8364
001b725c
6d8c744c
366417c3
126410c3
60376046
00ff131c
313c2954
554c01c7
408c0d00
0464325c
1004933c
60376186
600739c3
68cc1b54
002c245c
245c4d8f
4daf004c
006c245c
245c4dcf
4def008c
325c408c
68920464
0467325c
6d2c744c
402606c3
60063664
3f3c6037
2f5c1040
233c0001
735c805e
594c000e
06c3886c
23c318c3
46646066
c0764196
08040f56
bf96f016
71c350c3
802c7364
001b625c
6d8c704c
366416c3
126410c3
40374046
00ff131c
313c1454
514c01c7
6c8c6d00
0464335c
0100341c
40374186
704c68d2
05c36d2c
36644006
60376006
10403f3c
00012f5c
805e233c
000e635c
886c554c
17c305c3
606623c3
41964664
08040f56
0136f016
60c3bf96
736471c3
31cc802c
535c718c
a00703a1
64e91194
0e546027
0c546047
648d6869
44ed4046
704ca4ae
20266d4c
a0373664
61860073
3f3c6037
2f5c1040
233c0001
594c805e
06c3886c
23c317c3
46646026
80764196
08040f56
0136f016
50c3bf96
736471c3
31cc802c
635c718c
c00703a1
64e91494
11546027
0f546047
648d6869
64ad6889
64cd68a9
44ed4026
6d4c704c
366412c3
0073c037
60376186
10403f3c
00012f5c
805e233c
886c554c
17c305c3
602623c3
41964664
0f568076
00000804
bf967016
61c350c3
202c6364
658c45cc
03a1035c
60376186
0ff28006
40c368e9
02946047
606688ab
644c68ed
05c36d4c
36642006
00370006
10403f3c
00012f5c
805e233c
000e435c
886c554c
16c305c3
606623c3
41964664
08040e56
be96f016
52c360c3
736471c3
225c802c
4077001b
6d8c704c
366412c3
126410c3
60376046
00ff131c
313c3354
514c01c7
4c8c6d00
035c712c
30c30121
0020341c
21546007
0309025c
341c30c3
60070020
255c1a54
32c3002b
33647ca5
00e0331c
255c15b4
32c3003b
feb8321c
331c3364
0cb40700
6dac704c
25c306c3
30c33664
00b33264
40374346
62460073
0f5c6037
0f5c0001
2f5c0045
2f5c0021
794c004d
06c38c6c
2f3c17c3
60660080
42964664
08040f56
c0963016
4d2c602c
10003f3c
533ca006
ab0b805e
000e535c
535cab2b
414c001e
2fc3886c
466460a6
0c564096
00000804
bf967016
536451c3
2d2c602c
001b425c
fe50343c
331c3364
10b400e0
02be623c
321c36c3
3364feb8
0700331c
870e07b4
672e680b
c037c006
42460073
3f3c4037
6f5c1040
633c0001
414c805e
15c3886c
602623c3
41964664
08040e56
c0961016
10003f3c
233c4006
401c805e
435c00fb
201c000e
235c4290
435c001e
235c002e
414c003e
2fc3886c
46646126
08564096
00000804
bf96f016
42c350c3
636461c3
452c202c
37c3ebeb
001c341c
e037e186
13946007
0121725c
341c37c3
42260040
6bd24037
420c644c
143c6dcc
49490030
30c33664
60373264
10403f3c
00017f5c
805e733c
886c554c
16c305c3
602623c3
41964664
08040f56
bf96f016
61c350c3
802c6364
e7eb312c
341c37c3
e186001c
6007e037
715c1194
37c30121
0040341c
20372226
704c69d2
123c6dec
36640030
326430c3
3f3c6037
2f5c1040
233c0001
554c805e
05c3886c
23c316c3
46646026
0f564196
00000804
bf967016
61c350c3
202c6364
8beb452c
341c34c3
8186001c
6ff28037
0121425c
341c34c3
42260040
67d24037
6e0c644c
30c33664
60373264
10403f3c
00014f5c
805e433c
886c554c
16c305c3
602623c3
41964664
08040e56
bf967016
61c350c3
402c6364
135c692c
31c30121
0040341c
20372226
684c69d2
1f3c6e2c
36640050
326430c3
3f3c6037
2f5c1040
233c0001
554c805e
05c3886c
23c316c3
46646046
0e564196
00000804
bf967016
61c350c3
202c6364
435c652c
34c30121
0040341c
80378226
644c6bd2
123c6e4c
2f3c0030
36640050
326430c3
3f3c6037
2f5c1040
233c0001
554c805e
05c3886c
23c316c3
466460e6
0e564196
00000804
bf967016
61c350c3
202c6364
435c652c
34c30121
0040341c
80378226
644c6bd2
123c6e6c
2f3c0030
36640050
326430c3
3f3c6037
2f5c1040
233c0001
554c805e
05c3886c
23c316c3
466460e6
0e564196
00000804
bf96f016
61c350c3
802c6364
e7eb312c
341c37c3
e186001c
6007e037
715c1194
37c30121
0040341c
20372226
704c69d2
123c6e8c
36640030
326430c3
3f3c6037
2f5c1040
233c0001
554c805e
05c3886c
23c316c3
46646026
0f564196
00000804
bf967016
61c350c3
202c6364
435c652c
34c30121
0040341c
80378226
644c69d2
123c6eac
36640030
326430c3
3f3c6037
2f5c1040
233c0001
554c805e
05c3886c
23c316c3
46646026
0e564196
00000804
bd96f016
71c350c3
802c7364
001b625c
6d8c704c
366416c3
326430c3
40374046
40774006
331c40b7
0c5400ff
01c7333c
6d00514c
4e096c0c
6e294077
600660b7
3f3c6037
2f5c10c0
233c0001
635c805e
2f5c000e
2f5c0021
2f5c007d
2f5c0041
554c0085
05c3886c
23c317c3
466460a6
0f564396
00000804
bf967016
02c350c3
742c1364
40c34d2c
029e643c
341c36c3
64f20001
325c60c9
d009016d
341c36c3
6cf20002
0169325c
60e943c3
1a2c433c
4f5c8037
425c0001
3f3c016d
c0061040
805e633c
886c554c
23c305c3
46646026
0e564196
00000804
0136f016
70c3ba96
81c362c3
a02c8364
6d8c744c
001b125c
10c33664
60461264
131c6177
4c5400ff
01c7313c
6d00554c
8c8c6c8c
6ecc744c
26c307c3
30c33664
61773264
3c946007
123c26c3
31c3029e
0001341c
70096ff2
141c13c3
20b700f8
00413f5c
78c9700d
20b713a3
00411f5c
2809300d
341c31c3
60070002
50091094
341c32c3
60f700c7
00611f5c
58e9300d
19ac323c
3f5c6077
700d0021
323c5009
6ed20244
03f4323c
1f5c6137
300d0081
323c5909
603731ac
00013f5c
3f3c700d
1f5c1180
133c00a1
5d4c805e
07c3888c
23c318c3
46646026
80764696
08040f56
0136f016
60c3bf96
736471c3
31cc802c
535c718c
a00703a1
64e91394
10546027
0e546047
648d6869
64ed6046
6889a4ae
704c650d
20266d4c
a0373664
41860073
3f3c4037
2f5c1040
233c0001
594c805e
06c3886c
23c317c3
46646026
80764196
08040f56
0136f016
50c3bf96
736471c3
31cc802c
635c718c
c00703a1
64e91694
13546027
11546047
648d6869
64ad6889
64cd68a9
650d68c9
44ed4026
6d4c704c
366412c3
0073c037
60376186
10403f3c
00012f5c
805e233c
886c554c
17c305c3
602623c3
41964664
0f568076
00000804
c096f016
71c350c3
602c7364
10004f3c
243c4006
6d2c805e
00100f3c
01c0133c
b0bc4106
754c08cb
05c3cc6c
2fc317c3
66646126
0f564096
00000804
be967016
61c340c3
60066364
00053f5c
5f3c61ac
6c2c1000
15c30106
36644046
00100f3c
410615c3
08cbb0bc
ac6c714c
16c304c3
61262fc3
42965664
08040e56
0136f016
60c3bd96
836481c3
001b725c
10705f3c
200605c3
bebc40a6
982c0891
6d8c704c
17c306c3
30c33664
40463264
331c4037
175400ff
01c7333c
6d00514c
415c2c8c
88f202d1
28e505c3
b0bc40a6
803708cb
05c30113
40a62985
08cbb0bc
60376006
00012f5c
003d2f5c
00704f3c
000e745c
00a00f3c
10701f3c
b0bc40a6
794c08cb
06c3ac6c
24c318c3
56646106
80764396
08040f56
bf96f016
71c350c3
80067364
0030623c
542c02f3
01c7343c
6c80294c
033c6c8c
16c304c0
b0bc40a6
742c08cb
6d2c6c6c
366405c3
0010343c
4f5c6037
760c0001
34e46c29
3f3ce734
40061040
805e233c
886c554c
17c305c3
602623c3
41964664
08040f56
bd96f016
71c350c3
802c7364
cfeb712c
60376186
1194c007
10400f3c
0030123c
b0bc40e6
706c08cb
05c36d0c
08211f5c
10502f3c
c0373664
00013f5c
00253f5c
8c6c754c
17c305c3
00402f3c
46646026
0f564396
00000804
c0967016
42c350c3
636461c3
620c402c
313c2d09
294c01c7
0c2c6c80
64077049
34c30c94
019e133c
0275105c
143c0ae5
4c090040
08cbb0bc
10003f3c
233c4006
554c805e
05c3886c
2fc316c3
46646026
0e564096
00000804
bf967016
42c350c3
636461c3
620c402c
313c2d09
294c01c7
0c2c6c80
42467049
64074037
34c30d94
019e233c
03c542ad
0040143c
b0bc4c09
600608cb
3f3c6037
1f5c1040
133c0001
554c805e
05c3886c
23c316c3
46646026
0e564196
00000804
c096f016
71c350c3
4f3c7364
60061000
805e343c
6d2c602c
00100f3c
0240133c
b0bc4106
754c08cb
05c3cc6c
2fc317c3
66646126
0f564096
00000804
c0967016
61c340c3
60ac6364
04f0033c
0030123c
b0bc4106
2f3c08cb
60061000
805e323c
ac6c714c
16c304c3
60262fc3
40965664
08040e56
0736f016
70c3be96
a1c342c3
202ca364
3410a62c
cfeb652c
60776186
2c94c007
5489620c
0049835c
607760e6
243428e4
0040843c
6cac646c
019e143c
366428c3
326430c3
331cc077
169400ff
30097489
123c29c3
74893e9d
69806312
0010033c
82bc18c3
54890942
602532c3
1f5c6037
348d0001
3f3cc077
2f5c1080
233c0021
5d4c805e
07c3886c
23c31ac3
46646026
e0764296
08040f56
b896f016
42c350c3
736471c3
692c402c
20372186
20072da9
645c4194
684c002b
06c36d6c
366415c3
326430c3
60076037
345c3594
6132001b
08263f5c
088c363c
08363f5c
3f5c70e9
31e9084d
08451f5c
3f5c7109
0f3c0855
143c10b0
82bc0090
310b0942
08961f5c
3f5c712b
314b08a6
08b61f5c
3f5c716b
318b08c6
08d61f5c
3f5c71ab
742c08e6
6c6c6c6c
1f3c05c3
36641040
326430c3
1f5c6037
1f5c0001
754c0025
05c38c8c
2f3c17c3
60260040
48964664
08040f56
c0967016
61c340c3
602c6364
123c0d2c
82bc0030
2f3c0942
60061000
805e323c
ac6c714c
16c304c3
60262fc3
40965664
08040e56
be967016
61c350c3
602c6364
100c8e2c
6feb6d2c
41866037
6bf24077
2d29760c
9cbc2312
3f5c08cb
708d0001
40774017
10803f3c
00212f5c
805e233c
886c554c
16c305c3
602623c3
42964664
08040e56
0336f016
70c3fe96
836481c3
b94cc02c
68eb290b
23b431e4
31e4694b
383c2014
b58001c7
8d6c786c
35c32026
786c4664
1f5c2006
8cec0005
28c307c3
46646006
325c548c
60720404
0407325c
8bcb592c
602534c3
20066bce
00732077
40774246
00213f5c
029603c3
0f56c076
00000804
51c33016
802c5364
6c0c704c
366415c3
335c718c
604703a1
353c0854
514c01c7
6c0c6d00
4e8d4026
08040c56
ff963016
536451c3
6c6c602c
00052f5c
20468cec
600625c3
00064664
0c560196
00000804
fd96f016
e02c60c3
0373a006
01c7353c
6d005d4c
6e896c0c
602760b7
7c6c0d94
2f5c4006
8cec0005
3f5c06c3
13c30041
600625c3
353c4664
60770010
00215f5c
6c097a0c
e3b435e4
0f560396
00000804
fe96f016
51c362c3
602c5264
8c896e2c
40060c0c
02d34077
35e46009
20060b94
4c296080
23e478a2
20250594
f99420c7
60570213
e02573c3
2f5ce037
40770001
60570105
74e473c3
301ce814
607700ff
00217f5c
029607c3
08040f56
0136f016
80c3fd96
62c341c3
bd2ce02c
158d00c6
376e2006
574e5fe6
778e6366
0060053c
286c28c3
094282bc
728d6106
0c80001c
102f100f
0c80101c
03d6145c
508e4006
714d6006
0006716d
510e106f
40e634c3
095e233c
210603c3
0942a0bc
3f5c00b7
345c0041
0046025d
0265045c
326d2006
580d4026
386d382d
786e6406
188e0206
01e0043c
9cbc23e6
200608cb
7e0c32ad
23060c0c
08cb9cbc
00fb201c
301c570e
772e0848
0169355c
055c0006
341c0175
233c00c0
407703f5
00213f5c
016d355c
03d34006
32e46429
323c0c35
3d4c01c7
6c8c6c80
035c0006
200602d5
0407135c
01c7323c
6c001d4c
20066c0c
2e8d2e6d
0d4d0106
0010323c
2f5c6037
08c30001
6409220c
dfb432e4
80760396
08040f56
fd967016
326431c3
602c6077
940cae2c
20073489
6c6c2754
6f5c6cac
16c30021
30c33664
331c3264
1c5400ff
62c35489
c037dfe5
00011f5c
2f5c20b7
548d0041
1e1d643c
3f9d643c
51806312
631231c3
2c2c7180
7489282f
11806312
9cbc2106
039608cb
08040e56
60c37016
013351c3
f2bc05c3
798c0942
06c36c4c
366414c3
97f2942c
08040e56
42c31016
402c1364
01c7313c
6c80294c
2deb6c0c
4e8d4006
b8bc34c3
08560946
00000804
0736f016
60c3ff96
602c71c3
2e242d30
f52481c3
0070a73c
0473a026
353c582c
294c01c7
8c0c6c80
60277269
0ac30e94
0160143c
094288bc
326430c3
728966f2
60274166
02531294
47f25269
47eb19c3
341c32c3
69d20004
0010353c
536453c3
6c297a0c
dbb435e4
383c4006
62d24004
7a0cf324
21a66c29
35e42037
40373154
2e544167
353c582c
294c01c7
8c6c6c80
6c0c0c90
4e6d4026
306e3c0b
508e5c2b
306d3ca9
504d5c89
308d3cc9
0160033c
82bc1ac3
70490942
06946027
0400083c
82bc19c3
20260942
2dad39c3
6c6c782c
06c36d4c
25c317c3
40063664
3f5c4037
03c30001
e0760196
08040f56
fd96f016
326431c3
402c6037
2d09620c
01c7313c
6c80294c
ec0c8c2c
d04bb00b
43f24017
0413508e
13c36017
07942027
3f5c708e
345c0001
02d303bd
21c32017
07944087
708e6026
145c2046
019303bd
32c34017
604720c6
40170654
606732c3
20460394
35c3308e
0f5456e4
6c2c61ac
1f3c0046
20c300a0
0f5c3664
3aa00053
0a7c6ebc
33647400
345c6132
124903d6
094a0abc
00770264
00213f5c
025d345c
0261145c
4e27313c
333c4057
7dcf228d
0f560396
00000804
fe967016
32c340c3
32641364
402c6037
01c7313c
cc80294c
ac0c788c
4c09612c
341c32c3
60070002
60ac2854
0279135c
341c31c3
60070004
614c2054
1f3c6e6c
5fe60040
47c63664
2066400d
2f5c204d
406d0001
29eb580c
540b204e
342b406e
544b208e
40ae4332
402d4146
6c0c714c
205704c3
36644186
0e560296
00000804
fe963016
32c340c3
536451c3
60373264
4c09612c
341c32c3
60070002
60ac2054
0289235c
341c32c3
60070008
614c1854
1f3c6e6c
5fe60040
47c63664
4286400d
505c404d
2f5c001e
40ad0001
402d4086
6c0c714c
205704c3
366440c6
0c560296
00000804
ff967016
136440c3
313c402c
294c01c7
788ccc80
612caccc
32c34c09
0002341c
28546007
135c60ac
31c30279
0010341c
20546007
6e6c614c
5fe61fc3
47c63664
20a6400d
580c204d
105c29eb
540c001e
002f205c
105c342c
255c004f
205c0263
21a6006e
714c202d
04c36c0c
41e62017
01963664
08040e56
0136f016
50c3ff96
21c332c3
83c32364
602c8264
612c2d4c
34c38c09
0002341c
3e546007
435c60ac
34c30281
0040341c
36546007
01c7323c
708c8580
ec6ccc4c
6e6c614c
5fe61fc3
27c63664
40e6200d
700c404d
405c8deb
18c3001e
580b2ef2
002e205c
305c784b
9c0b003e
004e405c
105c3c4b
0193005e
205c4366
301c002e
305c0148
205c003e
305c004e
8166005e
754c802d
05c36c0c
41a62017
01963664
0f568076
00000804
fc963016
32c340c3
32641364
402c6037
01c7313c
4c80294c
612ca80c
31c32c09
0002341c
40546007
215c288c
323c0404
65d22004
699232c3
0407315c
235c70ac
32c30279
0040341c
2e546007
6e6c714c
1f3c04c3
5fe600c0
67c63664
2186600d
2f5c204d
406d0001
604e75eb
20773609
04352047
60cd6066
1f5c0093
20cd0021
a0b7b629
604735c3
20660435
009320ed
00412f5c
60c640ed
714c602d
04c36c0c
410620d7
04963664
08040c56
fe967016
32c360c3
236421c3
60373264
2d4c602c
8c09612c
341c34c3
60070002
60ac2c54
0279435c
341c34c3
60070008
323c2454
a58001c7
6e6c614c
00401f3c
36645fe6
47c640c3
6086400d
2f5c604d
406d0001
4deb740c
748c404e
133c00c5
41060610
08cbb0bc
702d6186
6c0c794c
205706c3
366441c6
0e560296
00000804
fb967016
63c350c3
20f71264
40b72264
01212f5c
3f5c4077
60370160
4c09612c
341c32c3
60070002
60ac3354
0281235c
341c32c3
60070008
614c2b54
1f3c6e6c
5fe60100
40c33664
600d67c6
404d4166
606d6026
00612f5c
3f5c408d
60ad0041
16c300c5
094282bc
00212f5c
043c518d
229700d0
094282bc
00013f5c
4246726d
754c502d
05c36c0c
42862117
05963664
08040e56
fa967016
63c350c3
21371264
40f72264
01411f5c
2f5c20b7
40770180
2c09612c
341c31c3
60070002
60ac3e54
0279235c
341c32c3
60070002
614c3654
1f3c6e6c
5fe60140
40c33664
600d67c6
204d2046
406d4026
00813f5c
1f5c608d
20ad0061
16c300c5
094282bc
00412f5c
41a6518d
6ad26097
00d0043c
409722d7
08cbb0bc
21c32097
3f5c41a5
71210021
323c4025
6037ffe0
00011f5c
754c302d
05c36c0c
36642157
0e560696
00000804
0336f016
70c3fd96
81c332c3
32648364
20306077
4d4c39c3
cc09612c
341c36c3
60070002
60ac6354
0279135c
341c31c3
60070001
383c5b54
c98001c7
6e6c614c
00801f3c
36645fe6
47c650c3
6026400d
1f5c604d
206d0021
6d097e0c
129438e4
c006782c
2026c04e
4d6920cd
010540ed
00c0133c
094282bc
d50ed4ee
6006d52e
580c04b3
186c988c
d44ec9eb
313c2aa9
7fe50b0d
f88c133c
3f5c2037
13c30001
c08934cd
053cd4ed
123c0080
82bc0160
700c0942
34ee2c0b
4c2b700c
700c550e
63326c4b
345c752e
768d0289
d42dc266
6c0c7d4c
209707c3
366442a6
26d218c3
698c29c3
635cc006
039603b6
0f56c076
00000804
41c31016
6b86442b
4107311c
3fe64c0e
311c6346
2c0e4107
6045508b
321c4c0e
2c0e0080
618650ab
4107311c
321c4c0e
2c0e008e
644650cb
4107311c
600c4c0e
335c6cac
321c09c4
611200b9
236423c3
311c6746
4c0e4107
4c0e6045
9880201c
4103211c
341c680b
680efffd
08040856
6006400b
4107311c
5fe64c0e
00a0321c
60854c0e
404b4c0e
009e301c
4107311c
406b4c0e
4c0e6085
00000804
fe961016
136432c3
213c3264
141c40cb
01000007
60266cd2
100d433c
20098077
807741a3
00212f5c
0173400d
31236026
203713e3
12834009
3f5c2037
600d0001
08560296
00000804
1364ff96
40cb213c
0074313c
313c2122
133c308d
20370014
00012f5c
019602c3
00000804
311c63c6
0c0b4107
2000041c
00000804
0180201c
4107211c
600e680b
604d680b
00000804
301cff96
311c9892
6c0b4103
0010361c
090b233c
3f5c4037
03c30001
08040196
0136f016
70c3fe96
000b53c3
7e0530c3
036403c3
63c36820
340f6364
0010303c
7ffe101c
f3ff111c
201c3183
211c8000
32a30c00
05c3744f
60776026
20570653
406721c3
60260494
0a336037
333c6132
9d8000c7
12c34057
0001141c
0010313c
3a1d243c
60570205
821c83c3
8f5c0001
44f20027
00370046
343c0753
400f159d
0010233c
7ffe101c
f3ff111c
101c2183
111c8000
21a30c00
79a0404f
636463c3
00213f5c
cc94c007
7e056412
684c5580
684f6e72
311c67c6
6c0b2100
0001341c
40374086
13946007
236425c3
0092301c
2100311c
253c4c0e
6045808c
67464c0e
2100311c
0081001c
c0370c0e
00011f5c
029601c3
0f568076
00000804
fd963016
51c342c3
20065264
005d1f5c
00593f5c
0010133c
2f5c2037
40770001
00211f5c
005d1f5c
f33563a7
0004f524
00040004
301c400b
311c020e
4c0e4107
6045402b
404b4c0e
4c0e6045
6045406b
408b4c0e
4c0e6045
604540ab
40cb4c0e
4c0e6045
604540eb
101c4c0e
111c0200
640b4107
fff0253c
ff00341c
41ac323c
ff00341c
640e6472
0202201c
4107211c
341c680b
7dd20002
021e301c
4107311c
700e6c0b
0220301c
4107311c
702e6c0b
0222301c
4107311c
704e6c0b
0224301c
4107311c
706e6c0b
0226301c
4107311c
708e6c0b
0228301c
4107311c
70ae6c0b
022a301c
4107311c
70ce6c0b
022c301c
4107311c
70ee6c0b
0004f324
00040004
0c560396
00000804
52c37016
601c5264
611c9884
980b4103
301c400b
311c9888
4c0e4103
6045402b
404b4c0e
4c0e6045
6045406b
42644c0e
422c313c
780e3364
311c6706
ac0e4107
08040e56
311c61c6
201c4107
4c0e009f
311c6186
201c4107
4c0e0240
201c6a05
4c0e0096
311c6386
201c4107
4c0ee19f
6c4b61ec
07546067
00a8301c
4107311c
4c0e4026
00000804
ff963016
416442c3
ac8c600c
311c6586
40064107
6dc54c0e
00c0201c
01c34c0e
094a84bc
60660364
03e46037
24c31e35
301c2364
311c80b2
4c0e4103
86a4201c
4103211c
3364680b
680e6372
311c6446
40264107
355c4c0e
641211c4
000f351c
11c7355c
60376006
00012f5c
019602c3
08040c56
ff96f016
736472c3
400c3364
a84cc88c
211c4586
680e4107
009a301c
4107311c
00c0201c
055c4c0e
84bc01c9
0364094a
1c350127
055c966c
6abc01c9
40e4094a
301c1554
311c0180
ec0e4107
311c6446
40264107
365c4c0e
641211c4
000f351c
11c7365c
60376006
40660073
3f5c4037
03c30001
0f560196
00000804
50c3f016
0271701c
08958ebc
6120550c
080c433c
0271601c
3470341d
f5b46127
101c0006
c2bc0138
141d094a
00063460
2d00548c
094aa8bc
08958ebc
6120552c
080c433c
3460341d
f7b46127
101c0026
c2bc0138
301c094a
141d0271
00263430
2d0054ac
094aa8bc
08040f56
40c31016
84bc0006
303c094a
3364ed10
f9b46247
08958ebc
0006110f
094a6abc
201c108f
211cffff
12c30fff
039401e4
508f4006
96bc0006
0364094a
002610cf
094a84bc
ed10303c
62473364
8ebcf9b4
112f0895
6abc0026
10af094a
ffff201c
0fff211c
01e412c3
40060394
002650af
094a96bc
10ef0364
08040856
41c31016
f0bc01c3
6006097c
4107311c
700e6c0b
311c6b86
6c0b4107
301c702e
311c009e
6c0b4107
301c704e
311c00a2
6c0b4107
6386706e
4107311c
708e6c0b
311c6186
6c0b4107
644670ae
4107311c
70ce6c0b
08040856
3f36f016
80c3f996
326432c3
25306137
1f5c2006
40d000dd
6c0c618c
01401f3c
c1573664
69ab29c3
a007aae9
60252494
78c37a8e
6c6b7ccc
6c000157
6157784f
0130233c
2c6b7ccc
79af6880
4c0d4046
5ac37ccc
ec6bb44b
133c77a0
09c3fec0
13e461ab
13c30235
0110313c
6006784e
04137aae
58c37a8e
6c6b74cc
6f80e157
6157784f
0140233c
0c6b74cc
79af6800
1ac374cc
4c6b244b
133c6520
59c3fec0
13e475ab
13c30235
0100313c
0006784e
41171aae
602732c3
52c31754
a04746d2
40671954
03932394
01c04f3c
00813f5c
ffde343c
a1174026
361c35c3
7fe50004
f88c033c
4f3c0433
ffe601c0
ffde743c
4f3cfe53
0aa601c0
ffde043c
4f3cfd93
5e0601c0
ffde243c
401cfcd3
411ca284
fc330013
b00979ac
9000ad21
0010323c
236423c3
37f23fe5
5dab79c3
044b1ac3
74cc58c3
60a02c6b
a0267d85
673523e4
64204285
a026e980
0140cf3c
30c30117
0004361c
b33c7fe5
07f3f88c
21772006
698c28c3
08c36c0c
36641cc3
604b0ac3
73e407c3
03c30235
088c353c
153c6037
333c0014
6c800037
0020d33c
3dc34157
3b9d263c
323c4017
6c800067
063c6045
df5c371d
003700a4
60776006
700901d3
40571dc3
4b846521
602532c3
60773364
32c34017
60377fe5
32f22017
353cfc20
60f70010
00615f5c
c194e007
253c0313
153c088c
323c0014
6c800067
e0066045
371d763c
0037323c
60456c80
063c0006
253c3b9d
40b70010
00415f5c
e835a0a7
d40f59c3
fc760796
08040f56
2264fe96
32644077
32c36037
05546027
32c34057
08946047
00012f5c
3f5c400d
640d0021
40060073
0296440d
00000804
326431c3
60272264
101c1a94
40873304
101c2b54
41473206
101c2754
41c72306
101c2354
41073302
101c1f54
41673106
101c1b54
41e71306
02d31894
15946007
40872206
101c1154
41470400
101c0d54
41670800
101c0954
41c74000
41e70554
101c0494
200e8000
6372600b
0804600e
4d8c600c
6025690c
0804690f
850c1016
24d2308c
6c2c618c
60063664
0856708f
00000804
4d4c600c
6025690c
0804690f
4d4c600c
6025690c
0804690f
fc967016
326431c3
a00c60f7
556c944c
21072809
760c0635
20a66e0c
05d33664
36c3c88b
688e6045
0010613c
1f5cc0b7
280d0041
6025728c
0002341c
19946007
0111245c
40074077
700c1694
16c3cc29
20372025
00012f5c
3f5c4c2d
720d0021
6e4c760c
5f5c2046
25c30061
00733664
d20dc026
145c2006
04960135
08040e56
fb96f016
a4ec200c
858c444c
6025710c
6a8c710f
0003341c
680c69f2
76c3cc29
e137e025
00816f5c
f029cc2d
e007e0f7
70093e94
2e356107
6e0c660c
366420c6
60277089
30ab1594
313c508b
23e4080c
313c0ff4
30ac100c
70af6c80
0379255c
40b74172
00413f5c
037d355c
70ab0213
d0ac6112
70af6f00
0379755c
041c07c3
007700fd
00211f5c
037d155c
50cd4006
733c0273
e0370010
00010f5c
2026100d
3f5c2a0d
325c0061
00d30135
ca0dc006
725ce026
05960135
08040f56
ff967016
41c362c3
13c34364
6bc61264
2100311c
533c6c0b
40860014
a0074037
80072c94
313c1b94
7e05200c
684c4180
684f6e72
236420c3
009e301c
2100311c
203c4c0e
6045808c
6b464c0e
2100311c
0881201c
80374c0e
313c0213
4180200c
301cc80f
43a38000
884f4364
0010313c
61806412
a037686f
00012f5c
019602c3
08040e56
240c31c3
2c2c200f
2c8b202f
0804208e
0136f016
70c3fe96
04f061c3
a50c852c
6c2c61ac
1fc30046
366420c3
304b502b
085421e4
601748a0
3320341d
704f6c80
504f0053
6c12704c
28c3704f
6d004bcc
7009704f
74af6c12
74cf6006
4bd25029
6c0c7d8c
1f3c07c3
36640040
748f6057
54cd5029
74ed6006
6e0c7a0c
202607c3
02963664
0f568076
00000804
0136f016
70c3fc96
