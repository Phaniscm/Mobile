002374dc
0444975c
0464875c
275c4026
7c6c1ea5
133c07c3
08bc0b40
60c30b54
64dc0007
501c0022
511c10f8
740c0000
001c8c0c
3d2c0098
301c4146
311c6318
46640017
00071d8f
002122dc
7daf6146
275c3d2c
e6bc4764
60c30b0e
84dc0007
375c0020
0c0c0764
01801f3c
6c4c5d8c
0abeb4bc
0ef25d8c
4cbc02c3
00070b1c
375c4074
b0c31ed2
4a1503e4
fe67601c
4bd23df3
8c4c740c
3d2c02c3
301c4146
311c6318
46640017
10f8301c
0000311c
8c0c6c0c
3d2c0a06
301c44a6
311c6318
46640017
00071d8f
001d22dc
7daf64a6
275c3d2c
5ebc4764
00070ace
475c1294
84f20764
fec3601c
3f3c3873
033c01c0
100cfe7e
5d8c13c3
a4bc704c
03d20ab1
36d360c3
72bc1d8c
20c30ace
1ee2375c
0200b01c
041523e4
fe66601c
21263533
201c21b7
275c0200
301c0587
311c10f8
6c0c0000
02c38c0c
44c63d2c
6318301c
0017311c
50c34664
0567075c
f2dc0007
a9c30018
9a3ca884
02860090
05c7075c
383c1c70
375c0c40
07c305a7
0b3ed2bc
000740c3
7c2c5254
0a89235c
440d19c3
00667dac
64a70177
40260354
0f5c4177
39c300a1
7c2c0c2d
0a89435c
16548087
04b48087
06948047
80a70113
80c71c54
801c2754
07130002
275c4286
7c6c05c7
00c4321c
05a7375c
640605d3
05c7375c
321c7c6c
375c00d8
801c05a7
401c0002
0473019e
075c0606
7c6c05c7
00f8321c
05a7375c
0002801c
019f401c
280602d3
05c7175c
321c7c6c
375c0128
801c05a7
401c0002
013301a0
183c05c3
44860b40
08cbb0bc
8b0684c3
61477dac
64861b94
0587375c
0200001c
07c31dcf
0b3ed2bc
075c0cd2
175c0564
275c05a4
34c305c4
0ab594bc
0587075c
19c30bc3
08bc1884
60460b3f
1ea5375c
64a77dac
275c1794
475c05a4
575c05c4
373c0564
60370b00
20773d8c
60b76006
613760f7
12c307c3
35c324c3
0b6d40bc
7dac60c3
1d946147
0764275c
0564175c
0584575c
01973ac3
483ccc00
373c0020
60370380
60777d8c
00b7080c
60f7684c
01370006
25c307c3
74bc7a00
60c30b7a
a4dcc007
2066000c
1ea5175c
61972ac3
7daca980
119464a7
0584b75c
28c30bc3
08bc3500
383c0b3f
15800020
0564175c
0584275c
08cbb0bc
901c7dac
61470000
301c2a94
311c10f8
6c0c0000
1dcc8c0c
44c63d2c
6318301c
0017311c
90c34664
92dc0007
383c0009
35800020
b0bc5dcc
7dcc08cb
0564475c
0584175c
5d8c2037
07c34077
23c319c3
bcbc34c3
50c30b71
6a940007
375c6086
4bc31ea5
0ac34884
0020143c
37c341e6
0b444abc
00b0643c
202607c3
0b3eeabc
000730c3
643c3954
b01c0060
b11c10f8
1bc30000
8c0c640c
3d2c06c3
301c44c6
311c6318
46640017
b06680c3
3e540007
00501a3c
b0bc26c3
c03708cb
407742c6
60b76026
00f70006
1ac307c3
0466201c
debc38c3
60c30b57
640c1bc3
08c38c4c
44c63d2c
6318301c
0017311c
56c34664
0a15c007
07c30373
26c31ac3
0b5004bc
000750c3
60a61394
1ea5375c
0464375c
375c6f00
375c0467
341c1e44
a0060008
07c365f2
0b44d6bc
09c350c3
301c0fd2
311c10f8
6c0c0000
09c38c4c
44c63d2c
6318301c
0017311c
20064664
05a7175c
05c7175c
7ebc07c3
00930b51
56c3d066
05c3feb3
f0760796
08040f56
60c37016
4f540007
165c0085
f2bc2584
063c0b43
165c1900
f2bc2584
065c0b43
0fd224c4
10f8301c
0000311c
8c4c6c0c
2584165c
301c40c6
311c66e4
46640017
4a40063c
0ba7e6bc
10f8401c
0000411c
ac4c700c
2464065c
2584165c
301c45a6
311c66e4
56640017
ac4c700c
2644065c
2584165c
301c4666
311c66e4
56640017
8c4c700c
26a4065c
2584165c
301c4666
311c66e4
46640017
2544065c
200604d2
0aa318bc
08040e56
60c37016
0b3f74bc
200606c3
0b54ecbc
7ebc06c3
365c0b51
341c1e44
60070040
18cc1254
0b1c08bc
10f8301c
0000311c
8c4c6c0c
392c18cc
301c4406
311c66bc
46640017
10f8401c
0000411c
ac4c700c
392c182c
301c43c6
311c66bc
56640017
ac4c700c
392c186c
301c45c6
311c66bc
56640017
8c4c700c
04e4065c
4206392c
66bc301c
0017311c
063c4664
101c2c00
b8bc0104
065c0b06
05d20704
0724165c
0b06b8bc
10f8501c
0000511c
8c4c740c
0704065c
41e6392c
66bc301c
0017311c
740c4664
065c8c4c
392c06c4
301c41e6
311c66bc
46640017
0639265c
365c47f2
341c1e24
60070010
501c1b54
511c10f8
740c0000
065c8c4c
392c0684
301c41e6
311c66bc
46640017
8c4c740c
0644065c
41e6392c
66bc301c
0017311c
60064664
4745365c
0abc06c3
065c0ba8
00071f44
e6bc1254
301c0b1c
311c10f8
6c0c0000
065c8c4c
392c1f44
301c4146
311c66bc
46640017
03e1265c
06c345d2
4abc2026
365c0b4e
64d204c1
b4bc06c3
065c0b44
365c1f24
30e41f04
7abc0354
065c0bad
7abc1f04
065c0bad
00071f84
365c1554
63d22011
0ad2b6bc
10f8301c
0000311c
8c4c6c0c
1f84065c
44a6392c
66bc301c
0017311c
065c4664
00071fa4
265c1554
43d22019
0ad2b6bc
10f8301c
0000311c
8c4c6c0c
1fa4065c
44a6392c
66bc301c
0017311c
065c4664
00071fc4
365c1554
63d22021
0ad2b6bc
10f8301c
0000311c
8c4c6c0c
1fc4065c
44a6392c
66bc301c
0017311c
065c4664
392c4784
0b92e4bc
4884065c
301c0cd2
311c1110
6c0c0000
07c4335c
40063664
4887265c
4080063c
0b823ebc
1371365c
1a546007
10f8301c
0000311c
8c4c6c0c
0b44065c
4726392c
66bc301c
0017311c
363c4664
365c16e0
40060b47
1375265c
365c6006
0e560b66
00000804
50c37016
10f8601c
0000611c
8c4c780c
35cc000c
301c4166
311c6718
46640017
0ad215ac
8c4c780c
43c635cc
6718301c
0017311c
601c4664
611c10f8
780c0000
14ec8c4c
41e635cc
6718301c
0017311c
780c4664
14ac8c4c
41e635cc
6718301c
0017311c
142c4664
08bc0dd2
780c0b1c
142c8c4c
440635cc
6718301c
0017311c
053c4664
e6bc02c0
053c0ba7
e6bc0240
053c0ba7
e6bc0280
158c0ba7
0ba794bc
0444055c
e4bc35cc
0e560b92
00000804
50c37016
0080603c
cabc06c3
09d20b23
331c748c
2294fe63
d4bc05c3
02130b83
433c746c
946ffff0
ccbc06c3
80070b23
05c31594
0b83d4bc
c8bc06c3
301c0b23
311c10f8
6c0c0000
05c38c4c
424635cc
670c301c
0017311c
0e564664
00000804
50c37016
000c61c3
2cbc03d2
05c30b84
0b8292bc
10f8301c
0000311c
8c4c6c0c
16c305c3
301c4226
311c669c
46640017
08040e56
ff967016
51c340c3
200662c3
0098201c
0891b0bc
4026b00f
91cf506f
01f4301c
245c730f
043c0265
c6bc0080
00070b23
301c0615
708ffe63
06d312c6
245c4806
301c0276
345c0080
43860286
0296245c
345c6406
201c0326
211c382c
52af0017
36bc301c
0017311c
b44972cf
35c3a037
0a946027
00012f5c
023d245c
345c32c3
245c0225
7fc60245
0427345c
b6bc06c3
30c30ba7
001c118f
66d2fe99
012c201c
04a7245c
01960006
08040e56
41c31016
34542087
0dd42087
1b542027
04d42027
11542007
204701d3
20671d54
04130a94
305420c7
287420c7
325420e7
36542107
07930006
672c101c
0017111c
06734026
6730101c
0017111c
b0bc4046
04c308cb
101c05b3
111c6734
40660017
101c0493
111c6738
40860017
101c03d3
111c6740
40a60017
101c0313
111c6748
40c60017
101c0253
111c6750
40e60017
101c0193
111c6758
41060017
101c00d3
111c6764
41260017
08cbb0bc
08560026
00000804
40c33016
ac2c604c
00d34006
20066500
038d135c
304c4025
f97425e4
2e2510cc
f6bc25c3
20c30b1b
013308d2
6d00704c
135c2006
4025038d
f97425e4
08040c56
60c3f016
305c71c3
a00615c9
10546047
15e9405c
02c0021c
b0bc24c3
063c08cb
3e003000
b0bc24c3
543c08cb
465c080c
063c1583
3e803400
b0bc24c3
b60008cb
3600063c
24c33e80
08cbb0bc
465cb600
063c1593
3e803800
b0bc24c3
760008cb
3900063c
24c33d80
08cbb0bc
15c9365c
07946047
3a00063c
41062006
0891b0bc
0f560006
00000804
3f36f016
80c3fd96
15e9105c
1583205c
105c6500
6c801593
61e56112
210c133c
501c2037
511c10f8
740c0000
02868c0c
44c62006
6784301c
0017311c
00774664
8c0c740c
20060886
301c44c6
311c6784
46640017
740c90c3
0f268c0c
44c62006
6784301c
0017311c
a0c34664
8c0c740c
0090001c
44c62006
6784301c
0017311c
00b74664
8c0c740c
20060b86
301c44c6
311c6784
46640017
740cc0c3
0c068c0c
44c62006
6784301c
0017311c
d0c34664
4bd24057
69d239c3
27d21ac3
45d24097
63d23cc3
66940007
2fd22057
10f8301c
0000311c
8c4c6c0c
200601c3
301c44c6
311c6784
46640017
4fd229c3
10f8301c
0000311c
8c4c6c0c
200609c3
301c44c6
311c6784
46640017
6fd23ac3
10f8301c
0000311c
8c4c6c0c
20060ac3
301c44c6
311c6784
46640017
2fd22097
10f8301c
0000311c
8c4c6c0c
200601c3
301c44c6
311c6784
46640017
4fd22cc3
10f8301c
0000311c
8c4c6c0c
20060cc3
301c44c6
311c6784
46640017
3dc3d066
62dc6007
301c000b
311c10f8
6c0c0000
0dc38c4c
44c62006
6784301c
0017311c
d0664664
0cc314b3
0b00eebc
ecbc0dc3
60c30b1d
55940007
644c18c3
133c09c3
46062710
08cbb0bc
bf5c7ac3
56c30044
0300693c
0ac307f3
ccbc15c3
e0250b84
3d540007
0010453c
684c28c3
133c07c3
46062710
08cbb0bc
644c18c3
0300073c
0300133c
b0bc4406
28c308cb
073c684c
133c0500
44060100
08cbb0bc
1ac30dc3
0710253c
0b1ddabc
20570dc3
0b1dcabc
205706c3
b0bc4286
0cc308cb
488619c3
0b05a6bc
1bc30cc3
0b055cbc
0010b21c
601754c3
51e413c3
0893bf74
fed2601c
10f8501c
0000511c
8c4c740c
20060057
301c44c6
311c6784
46640017
8c4c740c
200609c3
301c44c6
311c6784
46640017
8c4c740c
20060ac3
301c44c6
311c6784
46640017
8c4c740c
20060097
301c44c6
311c6784
46640017
8c4c740c
20060cc3
301c44c6
311c6784
46640017
8c4c740c
20060dc3
301c44c6
311c6784
46640017
08c300f3
46bc2097
60c30b85
06c3f753
fc760396
08040f56
3f36f016
90c3fa96
ac30604c
10f8501c
0000511c
8c0c740c
20060286
301c44c6
311c6770
46640017
740c00b7
001c8c0c
20060214
301c44c6
311c6770
46640017
740c80c3
001c8c0c
20060243
301c44c6
311c6770
46640017
740c70c3
0b868c0c
44c62006
6770301c
0017311c
a0c34664
8c0c740c
20060c06
301c44c6
311c6770
46640017
4097b0c3
38c348d2
e5d266d2
43d22ac3
55940007
6fd26097
10f8301c
0000311c
8c4c6c0c
20060097
301c44c6
311c6770
46640017
4fd228c3
10f8301c
0000311c
8c4c6c0c
200608c3
301c44c6
311c6770
46640017
301cefd2
311c10f8
6c0c0000
07c38c4c
44c62006
6770301c
0017311c
3ac34664
301c6fd2
311c10f8
6c0c0000
0ac38c4c
44c62006
6770301c
0017311c
d0664664
40072bc3
000bf2dc
10f8301c
0000311c
8c4c6c0c
20060bc3
301c44c6
311c6770
46640017
15d3d066
eebc0ac3
0bc30b00
0b1decbc
000760c3
29c36094
08c3684c
0710133c
b0bc2dc3
3d3c08cb
bd800010
0410cd3c
28c346c3
40772d84
01402d3c
0f3c4037
14c300f0
0b84ccbc
43540007
07c38025
00f01f3c
b0bc24c3
29c308cb
1e00684c
0710133c
b0bc2dc3
29c308cb
05c3684c
0100133c
b0bc4406
29c308cb
053c684c
133c0200
44060300
08cbb0bc
17c30bc3
dabc2cc3
0bc30b1d
cabc2097
00570b1d
42862097
08cbb0bc
18c30ac3
a6bc4017
29c30b05
6f00684c
133c0ac3
5cbc2710
a0250b05
0001c21c
8067c205
0873b994
fed2601c
10f8401c
0000411c
ac4c700c
20060097
301c44c6
311c6770
56640017
ac4c700c
200608c3
301c44c6
311c6770
56640017
ac4c700c
200607c3
301c44c6
311c6770
56640017
ac4c700c
20060ac3
301c44c6
311c6770
56640017
8c4c700c
20060bc3
301c44c6
311c6770
46640017
09c3c6f2
0b8526bc
015360c3
26bc09c3
00d30b85
8abc09c3
60c30b85
06c3f793
fc760696
08040f56
1e24305c
1000341c
fabc64d2
00730b9a
0b86fcbc
00000804
0f36f016
60c3ff96
72c351c3
bf5c83c3
af5c0144
935c0164
6d090003
53946027
16540007
6007600c
002644dc
10f8301c
0000311c
8c0c6c0c
0104001c
43e61ac3
6790301c
0017311c
180f4664
a0074a53
740c1654
24dc6007
301c0025
311c10f8
6c0c0000
001c8c0c
1ac30104
301c43e6
311c6790
46640017
4813140f
0001b31c
c7d20e94
173c180c
29c30800
0aa144bc
1354a007
173c140c
01930a00
180cc7d2
0a00173c
44bc29c3
a7d20aa1
173c140c
29c30800
0aa144bc
6026c3d2
a3d2798d
358d2026
690928c3
14dc6087
c0070008
782c1654
74dc6007
301c0021
311c10f8
6c0c0000
001c8c0c
1ac30190
301c43e6
311c6790
46640017
40b3182f
1654a007
6007742c
002054dc
10f8301c
0000311c
8c0c6c0c
0190001c
43e61ac3
6790301c
0017311c
142f4664
b31c3e73
25940001
1154c007
10fc301c
0000311c
8e4c6c0c
173c182c
273c0800
60060c00
00074664
002024dc
3554a007
10fc301c
0000311c
8e4c6c0c
173c142c
273c0a00
60260d00
00074664
3df32654
1154c007
10fc301c
0000311c
8e4c6c0c
173c182c
273c0a00
60060d00
00074664
001de4dc
1154a007
10fc301c
0000311c
8e4c6c0c
173c142c
273c0800
60260c00
00074664
001cc4dc
6026c3d2
a3d2798d
358d2026
690928c3
14dc60e7
c0070008
784c1654
d4dc6007
301c0019
311c10f8
6c0c0000
001c8c0c
1ac30130
301c43e6
311c6790
46640017
3173184f
1654a007
6007744c
0018b4dc
10f8301c
0000311c
8c0c6c0c
0130001c
43e61ac3
6790301c
0017311c
144f4664
b31c2f33
25940001
1154c007
18c3784c
2006440b
03c32037
0800173c
0c00373c
0b1e8cbc
600730c3
0017e4dc
3554a007
18c3744c
2026440b
03c32037
0a00173c
0d00373c
0b1e8cbc
600730c3
2d732654
1154c007
18c3784c
2006440b
03c32037
0a00173c
0d00373c
0b1e8cbc
600730c3
0015a4dc
1154a007
18c3744c
2026440b
03c32037
0800173c
0c00373c
0b1e8cbc
600730c3
001484dc
4026c3d2
a3d2598d
758d6026
650918c3
74dc6107
c0070008
784c1654
34dc6007
301c0012
311c10f8
6c0c0000
001c8c0c
1ac30130
301c43e6
311c6790
46640017
2233184f
1654a007
6007744c
001114dc
10f8301c
0000311c
8c0c6c0c
0130001c
43e61ac3
6790301c
0017311c
144f4664
b31c1ff3
27940001
1354c007
173c184c
38c30800
42bc4c0b
30c30b1e
f4dc6007
073c000f
173c0e80
40860c00
08cbb0bc
3954a007
173c144c
38c30a00
42bc4c0b
30c30b1e
b4dc6007
073c000e
173c0ec0
04d30d00
1354c007
173c184c
38c30a00
42bc4c0b
30c30b1e
94dc6007
073c000d
173c0e80
40860d00
08cbb0bc
1354a007
173c144c
38c30800
42bc4c0b
30c30b1e
54dc6007
073c000c
173c0ec0
40860c00
08cbb0bc
2026c3d2
a3d2398d
558d4026
650918c3
73946127
1654c007
6007784c
000a44dc
10f8301c
0000311c
8c0c6c0c
0130001c
43e61ac3
6790301c
0017311c
184f4664
a0071253
744c1654
24dc6007
301c0009
311c10f8
6c0c0000
001c8c0c
1ac30130
301c43e6
311c6790
46640017
1013144f
0001b31c
cfd21e94
173c184c
38c30800
0cbc4c0b
073c0a9a
173c0e80
40860c00
08cbb0bc
2b54a007
173c144c
38c30a00
0cbc4c0b
073c0a9a
173c0ec0
03930d00
184ccfd2
0a00173c
4c0b38c3
0a9a0cbc
0e80073c
0d00173c
b0bc4086
afd208cb
173c144c
38c30800
0cbc4c0b
073c0a9a
173c0ec0
40860c00
08cbb0bc
2026c3d2
a3d2398d
558d4026
6006c4d2
07a7375c
a00705c3
20063a54
0787175c
06b301c3
06731066
6007780c
ffdad4dc
740cff53
f4dc6007
feb3ffdb
6007782c
ffdfa4dc
742cfe13
c4dc6007
fd73ffe0
6007784c
ffe744dc
744cfcd3
64dc6007
fc33ffe8
6007784c
ffeee4dc
744cfb93
04dc6007
faf3fff0
6007784c
fff6d4dc
744cfa53
f4dc6007
f9b3fff7
f0760196
08040f56
fd963016
204740c3
20670a54
301c0c54
0885ff53
20274006
01131b94
0540203c
00930006
243c0885
345c0540
333c1e24
3264090b
712c6037
bfc66077
12c3a0b7
2c00243c
2b00343c
0b885abc
03c330c3
0c560396
00000804
ff961016
305c40c3
341c1e24
66d20010
0b49d8bc
b4dc0027
345c006b
331c1e59
52dc00cc
331c006b
84dc00c0
245c0048
40371e61
62dc44a7
2017000f
44a721c3
31c358b4
32dc2187
23c3001e
29b46187
40a712c3
002fa2dc
20a731c3
23c30db4
b2dc6067
12c30020
e5dc4067
2047002a
0068e4dc
401747b3
610732c3
001e02dc
410712c3
20e705b4
006824dc
40174293
612732c3
002822dc
94dc4147
56930067
13c36017
02dc2247
23c30018
11b46247
41c712c3
0015e2dc
21c731c3
0018b0dc
61e723c3
0024e2dc
14dc4227
32330066
13c36017
e2dc2287
23c30022
e0dc6287
12c30012
6f544467
14dc2487
1ad30065
32c34017
e2dc65c7
12c30036
20b445c7
252731c3
000802dc
652723c3
12c308b4
4a5444e7
65dc24e7
1e73000a
32c34017
a2dc6567
12c3002d
f0dc4567
31c3000c
82dc2587
65a7002e
0062a4dc
20176573
231c21c3
42dc00a0
31c3003b
00a0131c
23c311b4
72dc6607
12c3002a
60dc4607
31c30029
42dc2627
6647002e
006104dc
20175ed3
231c21c3
f2dc00ac
31c30034
00ac131c
331c06b4
14dc00a1
76730060
21c32017
00ae231c
003612dc
00af131c
005f64dc
40e66ef3
15c5245c
345c6026
208615cd
15d5145c
245c4106
345c15dd
021315e5
145c20e6
402615c5
15cd245c
345c6086
210615d5
15dd145c
245c4066
640615e5
15ed345c
145c2506
400615f5
15fd245c
345c6206
345c1586
345c1596
739315a6
145c20e6
402615c5
15cd245c
345c6086
210615d5
15dd145c
15e5245c
60e60213
15c5345c
145c2026
408615cd
15d5245c
345c6106
206615dd
15e5145c
245c4406
650615ed
15f5345c
145c2026
420615fd
1586245c
1596245c
15a6245c
60e66db3
15c5345c
145c2026
40a615cd
15d5245c
345c6106
145c15dd
260615e5
15ed145c
245c4506
600615f5
15fd345c
145c2406
42061586
60e6fc13
15c5345c
145c2026
40a615cd
15d5245c
345c6106
206615dd
15e5145c
245c4606
650615ed
15f5345c
02d32006
145c20e6
402615c5
15cd245c
345c60a6
210615d5
15dd145c
15e5245c
245c4606
650615ed
15f5345c
145c2026
440615fd
1586245c
efd36206
145c20e6
402615c5
15cd245c
345c60a6
210615d5
15dd145c
245c4066
660615e5
15ed345c
145c2506
402615f5
15fd245c
345c6406
22061586
40e61f13
15c5245c
345c6026
204615cd
15d5145c
245c4106
345c15dd
628615e5
15ed345c
145c2506
400615f5
15fd245c
345c6206
31331586
145c20e6
402615c5
15cd245c
345c6046
210615d5
15dd145c
15e5245c
245c4286
650615ed
15f5345c
145c2026
420615fd
1586245c
608629b3
15c5345c
145c2026
404615cd
15d5245c
345c6106
145c15dd
228615e5
15ed145c
245c4506
600615f5
60860d73
15c5345c
145c2026
404615cd
15d5245c
345c6106
145c15dd
0ab315e5
345c6026
200615c5
15cd145c
245c4046
610615d5
15dd345c
0c532026
145c2026
400615c5
15cd245c
345c6046
210615d5
15dd145c
245c4026
628615e5
15ed345c
145c2506
245c15f5
0ab315fd
145c2086
402615c5
15cd245c
345c6046
1f5c15d5
145c0001
406615dd
15e5245c
345c6286
250615ed
15f5145c
245c4006
630615fd
1586345c
18732017
245c4086
602615c5
15cd345c
145c2046
410615d5
15dd245c
00013f5c
15e5345c
145c2286
450615ed
15f5245c
345c6026
230615fd
1586145c
18d34106
345c6026
200615c5
15cd145c
245c4046
610615d5
15dd345c
145c2066
428615e5
15ed245c
345c6506
200615f5
15fd145c
245c4206
60061586
2026d0f3
15c5145c
245c4006
3f5c15cd
345c0001
210615d5
15dd145c
245c4066
628615e5
15ed345c
145c2506
402615f5
15fd245c
345c6206
20061586
1596145c
15a6145c
40e640b3
15c5245c
345c6026
204615cd
15d5145c
245c4106
345c15dd
3f5c15e5
345c0001
250615ed
15f5145c
02d34006
245c40e6
602615c5
15cd345c
145c2046
410615d5
15dd245c
15e5345c
345c6286
250615ed
15f5145c
245c4026
640615fd
1586345c
06732206
245c40e6
602615c5
15cd345c
145c2046
410615d5
15dd245c
345c6066
228615e5
15ed145c
245c4506
600615f5
40e602f3
15c5245c
345c6026
204615cd
15d5145c
245c4106
606615dd
15e5345c
145c2286
450615ed
15f5245c
345c6026
220615fd
1586145c
15a6145c
1596145c
40e63373
15c5245c
345c6026
204615cd
15d5145c
245c4106
606615dd
15e5345c
145c2286
450615ed
15f5245c
345c6006
240615fd
1586145c
245c4206
245c15a6
2f531596
345c60e6
202615c5
15cd145c
245c4046
610615d5
15dd345c
145c2066
428615e5
15ed245c
345c6506
202615f5
15fd145c
245c4406
62061586
15a6345c
1596345c
21062b33
15c5145c
245c4046
608615cd
15d5345c
15dd145c
19132026
145c2106
404615c5
15cd245c
345c60a6
145c15d5
202615dd
15e5145c
00012f5c
15ed245c
345c6506
200615f5
15fd145c
41060b53
15c5245c
345c6046
208615cd
15d5145c
15dd245c
245c4066
640615e5
15ed345c
145c2506
400615f5
41060bd3
15c5245c
345c6046
20a615cd
15d5145c
15dd245c
245c4066
660615e5
15ed345c
145c2506
400615f5
61060d13
15c5345c
145c2046
408615cd
15d5245c
15dd345c
345c6026
240615e5
15ed145c
245c4506
345c15f5
067315fd
245c4106
604615c5
15cd345c
145c20a6
245c15d5
402615dd
15e5245c
345c6606
250615ed
15f5145c
15fd245c
245c4406
62061586
41060373
15c5245c
345c6046
208615cd
15d5145c
15dd245c
245c4066
640615e5
15ed345c
145c2506
402615f5
15fd245c
345c6206
345c1586
208615a6
1596145c
410611f3
15c5245c
345c6046
20a615cd
15d5145c
15dd245c
245c4066
660615e5
15ed345c
145c2506
402615f5
15fd245c
345c6406
22061586
15a6145c
245c4086
145c1596
125315b6
345c6126
204615c5
15cd145c
245c4086
610615d5
15dd345c
145c2066
440615e5
15ed245c
345c6506
200615f5
15fd145c
245c4206
245c1586
608615a6
1596345c
21260df3
15c5145c
245c4046
608615cd
15d5345c
145c2106
406615dd
15e5245c
345c6406
250615ed
15f5145c
245c4006
620615fd
1586345c
612609b3
15c5345c
145c2046
408615cd
15d5245c
345c6106
206615dd
61260613
15c5345c
145c2046
408615cd
15d5245c
345c6026
345c15dd
240615e5
15ed145c
245c4506
600615f5
15fd345c
145c2206
145c1586
408615a6
1596245c
345c6106
049315b6
145c2126
404615c5
15cd245c
345c6086
202615d5
15dd145c
15e5145c
245c4406
650615ed
15f5345c
145c2006
440615fd
1586245c
345c6206
208615a6
1596145c
245c4106
345c15b6
331c1e59
d2dc00c0
331c0020
92dc00cc
345c0020
67271e61
001532dc
1eb46727
42dc62c7
62c70011
60a709b4
61473b54
60876d54
0020e4dc
66670993
001322dc
05b46667
54dc65e7
0f730020
72dc6687
66a7001c
001fe4dc
6d671393
001122dc
0bb46d67
42dc67a7
6ce7000b
000d02dc
f4dc6787
0ff3001e
009d331c
0014f2dc
009d331c
331c06b4
34dc009c
2493001e
009e331c
0015f2dc
009f331c
001da4dc
60262f73
15c5345c
145c2006
404615cd
15d5245c
15dd345c
15e5345c
345c6286
250615ed
15f5145c
245c4006
02b315fd
245c4026
600615c5
15cd345c
15d5245c
15dd245c
15e5245c
145c2206
460615ed
15f5245c
15fd345c
345c6206
20061586
1596145c
15a6145c
40863193
15c5245c
345c6026
204615cd
15d5145c
15dd345c
15e5345c
245c4286
650615ed
15f5345c
145c2006
430615fd
1586245c
0c536106
145c20e6
402615c5
15cd245c
345c6046
245c15d5
245c15dd
228615e5
15ed145c
245c4506
600615f5
15fd345c
145c2206
05331586
245c40e6
602615c5
15cd345c
145c2086
345c15d5
345c15dd
09b315e5
345c60e6
202615c5
15cd145c
245c4046
145c15d5
145c15dd
628615e5
15ed345c
145c2506
400615f5
15fd245c
345c6406
22061586
15a6145c
1596145c
40e62553
15c5245c
345c6026
208615cd
15d5145c
15dd345c
15e5345c
245c4406
650615ed
15f5345c
145c2006
440615fd
1586245c
345c6206
345c15a6
21731596
145c20e6
402615c5
15cd245c
345c6086
204615d5
15dd145c
15e5245c
245c4406
650615ed
15f5345c
145c2006
420615fd
1586245c
15a6245c
1596245c
60861d93
15c5345c
145c2026
404615cd
15d5245c
15dd245c
15e5145c
345c6286
250615ed
15f5145c
245c4006
630615fd
1586345c
f4732106
245c40e6
602615c5
15cd345c
145c2086
404615d5
15dd245c
15e5345c
f0f36406
245c40e6
602615c5
15cd345c
145c2046
145c15d5
345c15dd
428615e5
60e6f6f3
15c5345c
145c2026
404615cd
15d5245c
15dd245c
4106ed33
15c5245c
345c6046
208615cd
15d5145c
245c4026
245c15dd
640615e5
15ed345c
145c2506
400615f5
15fd245c
345c6206
345c1586
208615a6
1596145c
15b6345c
41061093
15c5245c
345c6046
20a615cd
15d5145c
245c4026
245c15dd
660615e5
15ed345c
145c2506
400615f5
15fd245c
345c6406
22061586
61060373
15c5345c
145c2046
408615cd
15d5245c
15dd145c
345c6026
240615e5
15ed145c
245c4506
600615f5
15fd345c
145c2206
145c1586
408615a6
1596245c
15b6145c
610608d3
15c5345c
145c2046
40a615cd
15d5245c
15dd145c
345c6026
260615e5
15ed145c
245c4506
600615f5
15fd345c
145c2406
42061586
15a6245c
345c6086
245c1596
047315b6
145c20e6
402615c5
15cd245c
345c6046
345c15d5
200615dd
15e5145c
245c4286
650615ed
15f5345c
15fd145c
145c2206
145c1586
145c15a6
345c1596
7e721e24
1e27345c
1561345c
18946067
1569245c
14544007
1e24345c
345c6c72
101c1e27
111c2e20
320f0017
08354027
345c6d72
00931e27
fe0c001c
00060053
08560196
00000804
01c330c3
023513e4
080403c3
ff967016
01c340c3
23c312c3
01536006
65c3a9a2
6503a5a2
6f5cc037
d1a10001
30e46025
0196f614
08040e56
402d4026
400d4066
00000804
402d4046
400d4066
00000804
602d6066
0804600d
0364fe96
20c30077
40374832
00012f5c
2f5c440d
442d0021
08040296
40291016
400942c3
422c323c
0856640e
00000804
00f7fc96
583220c3
2f5c40b7
440d0041
503240d7
2f5c4077
442d0021
483240d7
2f5c4037
444d0001
00612f5c
0496446d
00000804
28d220c3
1d84005c
0010303c
1d87325c
005c00f3
303c1da4
325c0010
08041da7
001c30c3
6007ff53
335c1354
002615d1
0e546047
05b46047
60270006
01130894
60870046
03c30554
025400a7
08041fe6
201c0364
211cff01
32c30000
029403e4
080407e6
50c37016
301c61c3
311c10f8
6c0c0000
02068c0c
456612c3
67a8301c
0017311c
07d24664
c02fa00f
610d6006
606f6006
08040e56
640d6009
08040026
02d230c3
03c3608b
00000804
60c3f016
000771c3
501c1854
511c10f8
740c0000
002c8c4c
301c4566
311c67b4
46640017
8c4c740c
17c306c3
301c4566
311c67b4
46640017
08040f56
006c0053
600c04d2
fc9431e4
00000804
4784005c
0b92d4bc
602603d2
0804610d
0136f016
61c350c3
10f8801c
0000811c
f46c0493
6027740c
64670454
01b31294
680c28c3
142c8c4c
456616c3
6798301c
0017311c
00b34664
16c3142c
0b92b6bc
680c28c3
05c38c4c
456616c3
6798301c
0017311c
57c34664
dc94a007
0f568076
00000804
40c37016
63c351c3
12c301c3
92bc23c3
20c30b92
40071066
300c1354
500f286f
0ed2086c
35e4600c
20c30354
606cff53
2006686f
16c3206f
0b92e4bc
0e560006
00000804
31c31016
201c42c3
09d2ff53
23c32466
16bc34c3
20c30b93
402602f2
085602c3
00000804
40c31016
4784005c
d4bc2466
00070b92
002c1354
10540007
101c600c
111cffff
21c30fff
089432e4
08f0301c
20061180
38bc512c
08560b93
00000804
0336f016
80c3fe96
72c331c3
60773264
33540007
60377fe5
00013f5c
2db46087
10f8901c
0000911c
680c29c3
00268c0c
456617c3
67e8301c
0017311c
60c34664
0007b066
3f5c1c54
600d0021
202608c3
37c326c3
0b9316bc
03f250c3
01f3a026
680c29c3
06c38c4c
456617c3
67e8301c
0017311c
00734664
ff53501c
029605c3
0f56c076
00000804
1f36f016
60c3fe96
92c3b1c3
80069264
0001c01c
58700753
44f229c3
60077909
b80c3354
88bc05c3
03640b92
188c303c
83848bc3
480928c3
303c4077
2c3c0074
4037300d
00017f5c
13c36057
1c5417e4
0040343c
436443c3
0454a027
0c94a467
343c0093
00d30010
19c3182c
0b92b0bc
43c36200
20574364
27a321c3
1f5c4077
38c30021
6ac32c0d
c694c007
029604c3
0f56f876
00000804
08040006
40c31016
42d201c3
000683f2
302c00d3
b0bc508b
108b08cb
08040856
0f36f016
60c3fe96
82c371c3
926493c3
b01ca006
0a130001
19c35870
590924f2
49544007
04c3980b
0b9288bc
203c0364
303c188c
1b3c0074
2077300d
4d2238c3
00213f5c
375423e4
3e8004c3
0b922ebc
0040353c
436443c3
6027780c
54c30554
0f946467
182c00d3
acbc3e00
00d30b92
3e00182c
fabc29c3
62000b93
536453c3
ffe0343c
3d801620
0b922ebc
88bc180b
03640b92
188c203c
0074303c
300d1b3c
38c32037
30c30d22
203713a3
00011f5c
212108c3
c0076ac3
05c3b094
f0760296
08040f56
0f36f016
a1c3b0c3
72c383c3
901c7364
911c10f8
29c30000
8c0c680c
18c30186
301c4566
311c67cc
46640017
000750c3
29c32254
8c0c680c
18c307c3
301c4566
311c67cc
46640017
142f60c3
29c30ef2
8c4c680c
18c305c3
301c4566
311c67cc
46640017
00f356c3
27c31ac3
08cbb0bc
7411f48e
f07605c3
08040f56
40c33016
236451c3
101c3264
4027feb8
54093d94
13544067
06b44067
09544027
1c944047
40870133
40a70f54
02331794
0200101c
201c0173
01b30400
0800001c
47a6045c
101c0273
145c1000
01d347a6
2000201c
47a6245c
04c30133
45e62046
0b59c0bc
fe82101c
13c30233
301c6fd2
118008f0
512c3409
0b9368bc
202710c3
04c30594
0b92dcbc
01c32006
08040c56
ff963016
236450c3
32644037
401c69f2
4007feb8
40266a94
4805205c
600c0593
0464335c
600743c3
60176054
25946007
08f0201c
13c30100
38bc552c
40c30b93
53940027
246605c3
0b92dcbc
1e44355c
0a1b343c
0a5b343c
1e47355c
1e24355c
323c4017
355c0a9b
744c1e27
00012f5c
0385235c
07338017
72bc4017
40c30b4b
355c0cf2
69721e44
1e47355c
1e24355c
355c6a72
05331e27
1e940047
08f0201c
20061500
38bc552c
40c30b93
1d940027
246605c3
0b92dcbc
1e44355c
0a1b343c
0a5b343c
1e47355c
1e24355c
0a9b343c
1e27355c
00270133
355c0894
303c1e44
355c0a9b
80061e47
019604c3
08040c56
3f36f016
70c3fe96
9f5c61c3
82c301a4
32648364
00076037
20077054
33c46e54
f88ca33c
64d23ac3
a00759c3
c93c6654
b93c0020
a0061300
df3c45c3
0b330040
662018c3
5cf46067
1f3c1a00
3cbc0060
343c0b92
43c30020
1a004364
3cbc1dc3
343c0b92
43c30020
2f5c4364
71000023
46d438e4
00333f5c
165461a7
0b546467
31946027
3a0007c3
00015f5c
a8bc35c3
01130b94
3a0007c3
00015f5c
f0bc35c3
50c30b94
1ac30433
1d542007
d2bc07c3
00070b3e
1a001854
3cbc1cc3
29c30b92
1f5c082b
31c30023
30e47fe5
240619f4
0b9202bc
343c20c3
0bc30020
b0bc3980
005308cb
1f5ca006
70800023
436443c3
48e4a9f2
00d3a614
ff53501c
501c0073
05c3feb8
fc760296
08040f56
40c31016
0cd230c3
0b3ec4bc
08f26026
1561345c
00fe331c
00260294
03c330c3
08040856
fe963016
51c340c3
0b95eebc
19540007
1754a007
60376006
045c6077
153c4784
2fc30020
0b9408bc
0020303c
436443c3
08358047
ffe0043c
2ebc15c3
00530b92
04c38006
0c560296
00000804
fe961016
600640c3
60776037
0b95eebc
6dd230c3
4784045c
40061fc3
0b93acbc
05d20364
0020303c
036403c3
08560296
00000804
fe967016
61c350c3
0b95eebc
60540007
5e54c007
00370006
05c30077
0b934abc
4784055c
0bd28046
0020163c
60262fc3
0b9408bc
0020303c
436443c3
0cd2140c
0444005c
3a0009d2
60262fc3
0b9408bc
43c36200
05c34364
0b3ed2bc
30540007
2c2b742c
2c542007
3a0001a6
0b922ebc
0020343c
436443c3
4c2b742c
004502c3
2ebc3a00
343c0b92
43c30020
742c4364
3a000c2b
0b922ebc
0020343c
436443c3
01534006
035c6500
1a210981
343c4025
43c30010
342c4364
23e4642b
8047f474
043c0835
16c3ffe0
0b922ebc
80060053
029604c3
08040e56
fe963016
eebc50c3
40c30b95
2e540007
60376006
05c36077
0b934abc
4784055c
07d240c3
40261fc3
0b93acbc
436440c3
0bd2140c
0444005c
1fc308d2
acbc4026
62000b93
436443c3
d2bc05c3
09d20b3e
0c2b742c
303c06d2
71800060
436443c3
343c85d2
43c30020
04c34364
0c560296
00000804
ff967016
41c350c3
603762c3
24f202d2
ff53001c
01c303b3
41a62006
0891b0bc
215705c3
0b9260bc
0040143c
0b9246bc
00013f5c
355c710d
712d1561
1569355c
06c3714d
00b0143c
0b922ebc
01960006
08040e56
0736f016
fdd8f21c
a1c350c3
73c392c3
12646f5c
ff53301c
32540007
21b08f3c
18c3c037
3f5c27c3
e6bc1244
05c30b96
0b9270bc
05c340c3
14bc16c3
30c30ba0
00406f3c
14c306c3
355c23c3
26bc15e9
30c30b1d
14940007
18c306c3
14bc41a6
30c30b1d
06c30df2
27c319c3
0b1d14bc
06f230c3
1ac306c3
0b1d04bc
03c330c3
0228f21c
0f56e076
00000804
40c37016
62c351c3
3a540007
38542007
36544007
65e7680c
606c3335
1c80033c
0b2566bc
033c706c
153c1680
4ebc0100
04c30b25
0b3ed2bc
00074486
345c1e54
608715d1
44860435
0a946107
033c706c
15c32240
0b2500bc
14940007
345c4406
60a715d1
706c0a94
2900033c
50bc15c3
30c30b24
66f24606
0006580f
001c0073
0e56ff53
00000804
3f36f016
0077fd96
b2c3a1c3
c4176037
10f8401c
0000411c
ac0c700c
20060606
301c44c6
311c6854
56640017
700c80c3
0606ac0c
44c62006
6854301c
0017311c
90c35664
8c0c700c
0214001c
44c62006
6854301c
0017311c
70c34664
45d228c3
63d239c3
35940007
4fd228c3
10f8301c
0000311c
8c4c6c0c
200608c3
301c44c6
311c6854
46640017
6fd239c3
10f8301c
0000311c
8c4c6c0c
200609c3
301c44c6
311c6854
46640017
e007d066
000b82dc
10f8301c
0000311c
8c4c6c0c
200607c3
301c44c6
311c6854
46640017
14f3d066
0754c087
c0a78606
c0270c54
00930894
8406c046
c00600d3
00738206
8286c026
ca40141d
da40341d
7f323dc4
2c3cc384
40b7fff0
16c307c3
60172bc3
0b1d26bc
000760c3
07c35594
43d72397
0b1d14bc
000760c3
07c34d94
04bc18c3
b0c30b1d
45940007
5bc3abc3
07c30813
24c318c3
0b1d14bc
000760c3
07c33b94
43d72397
0b1d14bc
000760c3
07c33394
04bc19c3
60c30b1d
2c940007
23c36097
0f94a2e4
6dd23dc3
26060dc3
0b9202bc
405730c3
19c30a80
b0bc23c3
02b308cb
0e806057
24c319c3
08cbb0bc
18c307c3
14bc24c3
60c30b1d
07c30df2
04bc18c3
60c30b1d
b60007f2
0001a21c
c014ace4
08c36bc3
b8bc2606
09c30b06
b8bc2606
07c30b06
0214101c
0b06b8bc
10f8401c
0000411c
ac4c700c
200608c3
301c44c6
311c6854
56640017
ac4c700c
200609c3
301c44c6
311c6854
56640017
8c4c700c
200607c3
301c44c6
311c6854
46640017
039606c3
0f56fc76
00000804
3f36f016
0177f996
4137d1c3
c4d760f7
a33c6025
a31c088c
75dc0100
45570012
41b74b00
0080231c
001205dc
00e0131c
0011c5dc
10f8501c
0000511c
8c0c740c
0100001c
44c62006
685c301c
0017311c
b0c34664
8c0c740c
0100001c
44c62006
685c301c
0017311c
c0c34664
8c0c740c
0080001c
44c62006
685c301c
0017311c
70c34664
8c0c740c
00e0001c
44c62006
685c301c
0017311c
80c34664
8c0c740c
00e0001c
44c62006
685c301c
0017311c
90c34664
68d23bc3
46d22cc3
38c3e5d2
000763d2
2bc35594
301c4fd2
311c10f8
6c0c0000
0bc38c4c
44c62006
685c301c
0017311c
3cc34664
301c6fd2
311c10f8
6c0c0000
0cc38c4c
44c62006
685c301c
0017311c
efd24664
10f8301c
0000311c
8c4c6c0c
200607c3
301c44c6
311c685c
46640017
4fd228c3
10f8301c
0000311c
8c4c6c0c
200608c3
301c44c6
311c685c
46640017
39c3d066
12dc6007
301c0009
311c10f8
6c0c0000
09c38c4c
44c62006
685c301c
0017311c
d0664664
08c31013
2dc32006
0891b0bc
200609c3
b0bc2dc3
0bc30891
2ac32117
08cbb0bc
32c340d7
0001341c
69a02ac3
41170cc3
2ac32980
08cbb0bc
249707c3
b0bc26c3
1f0008cb
45572517
08cbb0bc
6197e037
40266077
08c340b7
2bc31dc3
9abc3ac3
60c30b97
14940007
6197e037
40466077
09c340b7
2cc31dc3
9abc3ac3
60c30b97
015707f2
28c31dc3
08bc39c3
401c0b92
411c10f8
700c0000
0bc3ac4c
44c62006
685c301c
0017311c
700c5664
0cc3ac4c
44c62006
685c301c
0017311c
700c5664
07c3ac4c
44c62006
685c301c
0017311c
700c5664
08c3ac4c
44c62006
685c301c
0017311c
700c5664
09c38c4c
44c62006
685c301c
0017311c
00734664
ff7c601c
079606c3
0f56fc76
00000804
3f36f016
d0c3f996
417721b7
bf5c6137
8f5c0244
cf5c0264
9f5c0284
e5d702a4
80078597
a9c34454
501ca884
a31cff7c
48b40080
10f8301c
0000311c
8c0c6c0c
0080001c
44c62006
6850301c
0017311c
60c34664
0007b066
1bc33554
b0bc28c3
38c308cb
1cc31980
b0bc29c3
e06708cb
e10703f4
e0860294
af5cc037
e0b70027
21970dc3
61174157
0b979abc
301c50c3
311c10f8
6c0c0000
06c38c4c
44c62006
6850301c
0017311c
01934664
0007bf5c
00278f5c
0047cf5c
00679f5c
0b98aebc
05c350c3
fc760796
08040f56
0136f016
50c3ea96
72c361c3
4f3c83c3
04c30180
44062717
08cbb0bc
03800f3c
44062757
08cbb0bc
67fc301c
0017311c
61a66037
80b76077
60f76806
61376797
617767d7
16c305c3
38c327c3
0b99eabc
80761696
08040f56
0136f016
50c3ea96
72c361c3
4f3c83c3
04c30180
44062717
08cbb0bc
03800f3c
44062757
08cbb0bc
681c301c
0017311c
61a66037
80b76077
60f76806
61376797
617767d7
16c305c3
38c327c3
0b99eabc
80761696
08040f56
0736f016
60c3fc96
15e9a05c
1583905c
1593805c
10f8301c
0000311c
8c0c6c0c
00e0001c
44c62006
680c301c
0017311c
70c34664
0007b066
984c3054
d2bc06c3
39c30b3e
18c33a84
343c4c80
60370300
0100343c
00b76077
15d1365c
07c360f7
080c123c
2710243c
7cbc6606
50c30b9a
06c306f2
46bc17c3
50c30b85
10f8301c
0000311c
8c4c6c0c
200607c3
301c44c6
311c680c
46640017
049605c3
0f56e076
00000804
fc967016
804c60c3
d2bcb02c
343c0b3e
60370100
0300343c
00b76077
15d1365c
043c60f7
26062710
0710243c
50bc35c3
04f20b9a
a8bc06c3
04960b9a
08040e56
0136f016
70c3ed96
42c381c3
64b76606
01801f3c
04802f3c
0b9756bc
2c740007
101c04c3
111c682c
40860017
08922abc
06d20164
6840601c
0017611c
601c00b3
611c6830
7c4c0017
2710533c
07c38497
0b3ed2bc
61e6c037
3f3c6077
60b70180
013780f7
15d1775c
08c3e177
25c32186
eabc6606
13960b99
0f568076
00000804
080422af
080422cf
3f36f016
b1c3fb96
73c382c3
a2dc6007
0c0c000a
62dc0007
2289000a
22a921c3
412c313c
323c42c9
22e981ac
c1ac213c
d01c40f7
40870038
d01c0354
eebc004c
30c309f8
61373264
216713c3
301c0894
311c1118
6c0c0000
36646c8c
035c7c0c
10c30161
0169035c
40ac203c
0171135c
812c213c
0179035c
c12c903c
c01c68c3
89e40001
98c304b4
c6c3c006
323c4117
60b703c7
1110a01c
0000a11c
600c0ac3
1f5c2026
40060006
00252f5c
00068e6c
29c31bc3
46643dc3
000740c3
3cc35354
16546007
b98469a4
035c7c0c
10c30161
0169035c
40ac203c
0171135c
812c213c
0179035c
c12c303c
023463e4
2ac396c3
6e0c680c
20c604c3
366440d7
000750c3
3ac31754
680c4c0c
00976c2c
2e4b6c00
1c942007
1c0c6aac
366415c3
16540007
15c31c0c
12bc5c4c
00070a5e
301c1854
311c0ef0
4c0c0000
0bb4301c
0000311c
143c0c0c
26640040
2ac301b3
8fac680c
00811f5c
15c301c3
46644c0c
9f94c007
801c0073
08c3ffff
fc760596
08040f56
0f36f016
b0c3fe96
82c3a1c3
200643c3
0c0c2077
09f8eebc
926490c3
1118301c
0000311c
6c0c6c0c
535ca006
100c0125
f2dc0007
706c0009
4f946007
00401f3c
5cbc504c
20c30a5b
1fc606d2
14dc4027
12130009
2ccc6057
533c308f
f42bfa80
635c7780
155c002b
20c30293
323c0173
7580180c
0380eccb
0010723c
2f5ce037
32c30001
31e43364
60e4f314
032002b4
1110301c
0000311c
335c6c0c
366407a4
106f10c3
0bb4701c
0000711c
1c0c0ef2
1abc15c3
301c08e7
311c0b84
6c0c0000
222b001c
0ab33664
26c305c3
0a006abc
15c31c0c
08e71abc
51c3306c
47542007
708c102c
a006cc20
1bf485e4
ae89700c
aea975c3
43ac253c
273ceec9
aee9812c
c12c353c
608746c6
49460254
86e458c3
56c30235
0ac36800
25c32580
08cbb0bc
6e80702c
56e4702f
301c0f94
311c1110
6c0c0000
07c4335c
3664106c
306f2006
302f308f
2bc30293
1e79325c
0f356127
2dd219c3
000b931c
301c0a54
311c1118
6c0c0000
e0266c0c
0125735c
005305c3
02961fe6
0f56f076
00000804
0136f016
a16c61c3
10f8801c
0000811c
f40c0353
0bd2178c
680c28c3
16c38c4c
301c4366
311c68b4
46640017
680c28c3
05c38c4c
436616c3
68b4301c
0017311c
57c34664
e694a007
0f568076
00000804
07d230c3
fe98001c
03546027
fe92001c
00000804
40c33016
268651c3
0b06b8bc
0040043c
428615c3
08cbb0bc
0180043c
0140153c
b0bc4286
000608cb
08040c56
0136f016
71c360c3
400652c3
803c540f
08c30080
0b23cabc
000732c6
782c3e94
473c740f
02530140
17c30085
eabc4286
09f208cb
033c740c
14c30180
eabc4286
07d208cb
4c0c740c
140c540f
ed940007
6007740c
301c1a94
311c10f8
6c0c0000
8c0c580c
296c0686
301c4386
311c6878
46640017
09d2140f
06bc17c3
740c0b9d
4c0f582c
782f740c
ccbc08c3
740c0b23
63f22006
fed1101c
807601c3
08040f56
0336f016
42c361c3
8f5c53c3
200600e4
903c2c0f
09c30080
0b23cabc
0007f2c6
516c5a94
412c01b3
13c3796c
069421e4
394c0085
08cbeabc
740c06d2
540f4c0c
12f2140c
66d238c3
64d2740c
60076f8c
740c3d54
3a546007
02c0033c
0361135c
febc4006
00070aba
740c3154
0261135c
2c542007
04c0033c
0369135c
febc4026
00070aba
d40c2354
fcbc194c
70c30b9c
400728c3
301c1d54
311c10f8
6c0c0000
1bac8c0c
44c62006
6888301c
0017311c
18c34664
0cd2040f
4fac740c
740c442f
4fac2f8c
08cbb0bc
701c0073
09c3fe69
0b23ccbc
c07607c3
08040f56
3f36f016
90c3fb96
72c3d1c3
21372006
20b720f7
280f43d2
09c3282f
2f3c1dc3
1cbc0100
40c30b9d
24dc0007
e0370018
1dc309c3
3f3c4117
6cbc00c0
60c30b9d
fe69031c
001794dc
0c0c39c3
02c9105c
a1cc2fd2
e2dca007
54090016
a2dc4007
05c30016
08920ebc
c364c0c3
1dc30193
2cc385b0
c2dc4007
058c0015
82dc0007
50c30015
10f8101c
0000111c
19c3640c
8c0c440c
0800001c
4586296c
6864301c
0017311c
b0c34664
fed1601c
42dc0007
201c0014
211c10f8
680c0000
0f068c0c
44c62006
6864301c
0017311c
a0c34664
10f8101c
0000111c
8c0c640c
20060c06
301c44c6
311c6864
46640017
2ac380c3
000743d2
3ac33194
301c6fd2
311c10f8
6c0c0000
0ac38c4c
44c62006
6864301c
0017311c
18c34664
301c2fd2
311c10f8
6c0c0000
08c38c4c
44c62006
6864301c
0017311c
301c4664
311c10f8
6c0c0000
0bc38c4c
45862006
6864301c
0017311c
d0664664
0dc31e33
201c1bc3
02bc0800
29c30ab5
8e4c680c
f2dc8007
4dec000b
3f3c0037
60770080
15c302c3
3bc32cc3
50c34664
13dc0007
6097000b
d2dc6007
0ac3000a
4f062006
0891b0bc
1ac308c3
35c34097
0ab088bc
640c19c3
13c308c3
34bc4d6c
28c30ac4
6007680c
000964dc
18c30dc3
0aa7f8bc
f4dc0007
e0070008
101c1854
111c10f8
640c0000
440c19c3
05c38c0c
44c6296c
6864301c
0017311c
1c0f4664
bc2f06d2
25c32097
08cbb0bc
6a6c28c3
b93c8d50
0bc30080
0b23cabc
0007d2c6
00d76c94
19540007
0007038c
301c1054
311c10f8
6c0c0000
440c19c3
296c8c4c
301c4366
311c6864
46640017
1ac300d7
b0bc4f06
047308cb
10f8301c
0000311c
19c36c0c
8c0c440c
296c0f06
301c4366
311c6864
46640017
000700f7
1ac31054
b0bc4f06
40d708cb
2d6c6117
6117280f
4d6f40d7
698c4117
698f6025
a007a0d7
e0072254
7c0c2054
1d546007
10f8301c
0000311c
19c36c0c
8c0c440c
296c1c2c
301c4366
311c6864
46640017
40d7178f
69d26b8c
6baf7c2c
0f8c60d7
5c2c3c0c
08cbb0bc
fcbc0cc3
60c30b9c
ccbc0bc3
00730b23
fe91601c
10f8501c
0000511c
8c4c740c
20060ac3
301c44c6
311c6864
46640017
8c4c740c
200608c3
301c44c6
311c6864
46640017
2cd22097
080c29c3
68d2626c
366401ec
64c300b3
601c0073
06c3fe93
fc760596
08040f56
0336f016
81c370c3
301c92c3
311c10f8
6c0c0000
0a068c0c
44c62006
6898301c
0017311c
60c34664
0007b066
7c0c2254
235c18c3
6d6c02c1
0ab00cbc
fe91501c
07c30af2
29c316c3
0b9ddabc
06c350c3
0aa7a4bc
10f8301c
0000311c
8c4c6c0c
200606c3
301c44c6
311c6898
46640017
c07605c3
08040f56
0336f016
81c370c3
901cc02c
911c10f8
02930000
7c0cb80c
2d6c06c3
0b9cd4bc
680c29c3
8c4c5c0c
296c06c3
301c4386
311c68a8
46640017
c00765c3
073cec94
c8bc0080
38c30b23
10546007
10f8301c
0000311c
5c0c6c0c
07c38c4c
4586296c
68a8301c
0017311c
c0764664
08040f56
01c330c3
023513e4
080403c3
02d230c3
03c360cc
00000804
31c320c3
30e40006
001c15d4
4007ff53
025c1154
031c1404
0394febd
01530046
feb9031c
00660394
031c00b3
0294fea9
080400c6
4ed220c3
1e24325c
0010341c
23d262d2
24d265f2
2c00023c
023c0073
08043000
0336f016
91c370c3
83c362c3
ff53301c
31540007
4087a026
40871354
a04607d4
a2c64fd2
0b944067
a4a60173
08544127
414752c3
a2a60554
02544107
301ca066
311c10f8
6c0c0000
093c8c0c
18c30140
301c25c3
311c6a18
46640017
301c1c0f
09d2fed1
a08fc06f
303c0031
600f0140
60062051
c07603c3
08040f56
006930c3
0c0910c3
c0ac203c
213c2c29
2c49812c
412c013c
00000804
0ba062bc
341d6166
08040030
1e24305c
0b8b033c
00000804
08040006
28a4205c
0408021c
02c342f2
00000804
03c0303c
30c302f2
080403c3
68c4001c
0017011c
00000804
0ba086bc
0ba08cbc
00000804
0b5690bc
00000804
50c33016
16540007
25a1305c
12546007
0b823ebc
10f8301c
0000311c
8c4c6c0c
155c05c3
45462584
695c301c
0017311c
0c564664
00000804
3f36f016
50c3fa96
407761c3
901c6037
911c10f8
19c30000
8c0c640c
20060b86
301c44c6
311c6970
46640017
000780c3
000d02dc
0b00eebc
101c06c3
111c68cc
40660017
08922abc
616460c3
14dcc007
05c3000c
1498301c
0000311c
40e62c0c
08922abc
e1060164
0007b7c3
05c34554
149c301c
0000311c
41862c0c
08922abc
e3060164
38540007
301c05c3
311c1480
2c0c0000
2abc4166
01640892
b7c3e206
2a540007
301c05c3
311c1484
2c0c0000
2abc4166
01640892
b01ce306
00070010
05c31b54
1488301c
0000311c
41662c0c
08922abc
e4060164
0010b01c
29c30dd2
8c4c680c
16c308c3
301c44c6
311c6970
46640017
a7c30df3
c0069bc3
d784dbc3
0080cf3c
c6d20a93
1cc308c3
a6bc4206
08c30b05
44572017
0b05a6bc
25d22057
410608c3
0b05a6bc
1cc308c3
0b055cbc
01738026
1cc308c3
a6bc4206
08c30b05
5cbc1cc3
80250b05
32c34497
f37443e4
1ac38206
12542007
22060ac3
0b9feebc
2ac340c3
24d77d20
1cc30580
b0bc24c3
da0008cb
4206a4a4
39c38a20
17546007
15548007
14c309c3
0b9feebc
251750c3
3bc32cd2
220639a4
25174620
3cc30580
25c32d00
08cbb0bc
95a4da80
ac746de4
10f8301c
0000311c
8c4c6c0c
200608c3
301c44c6
311c6970
46640017
02546de4
06c3c006
fc760696
08040f56
ff961016
205c40c3
47321e41
1e24305c
0010341c
34dc6007
40070012
305c1094
68d20744
66d26c0c
0764305c
6c0c63d2
201c66f2
245cfec3
22331407
0464345c
15546007
d6bc04c3
045c0b44
00071407
001064dc
14c4345c
345c6af2
23c31e99
40374025
00013f5c
1e9d345c
1e99345c
745460c7
10b460c7
35546047
07b46047
27546007
b4dc6027
0553000e
46546087
54b46087
61470673
000a52dc
07b46147
7d546107
f5dc6107
0d530008
e2dc6187
6187000a
000a10dc
14dc61a7
1753000d
7ebc04c3
045c0b78
00071407
000c83dc
1e71345c
f53560c7
345c6026
40461e9d
1e9d245c
cebc04c3
045c0b51
00071407
000b64dc
345c6066
345c1e9d
341c1e24
69f20400
4cbc04c3
045c0b5b
00071407
000a64dc
245c4086
345c1e9d
341c1e24
69f20400
98bc04c3
045c0b49
00071407
000964dc
345c60a6
345c1e9d
341c1e24
69f20400
8abc04c3
045c0b7a
00071407
000864dc
245c40c6
245c1e9d
323c1e24
6bf24004
0204323c
04c368d2
0b50b2bc
1407045c
73940007
345c60e6
345c1e9d
341c1e24
68f20400
88bc04c3
045c0b50
00071407
41066494
1e9d245c
1e24345c
0400341c
019369d2
7ebc04c3
045c0b78
00071407
345c5474
61071e71
6126f635
1e9d345c
1e44345c
0100341c
04c368d2
0b5038bc
1407045c
41940007
245c4146
04c31e9d
0b5d6abc
1407045c
37940007
345c6166
04c31e9d
0b5cfcbc
1407045c
2d940007
245c4186
345c1e9d
341c1e24
69f20400
04c30193
0b787ebc
1407045c
1d740007
1e71345c
f6356107
345c61a6
714c1e9d
04c369d2
3664316c
04150007
1407045c
345c0193
341c1e24
00264000
04c367f2
0b687cbc
00530026
01961fe6
08040856
ff963016
305c40c3
341c1e24
60070010
000de2dc
0464305c
14546007
0b44d6bc
1407045c
34dc0007
345c000d
6af214c4
1e91245c
602532c3
2f5c6037
245c0001
345c1e95
60a71e91
60a76e54
604711b4
60474f54
600707b4
60271d54
000b84dc
60670493
60874e54
000b24dc
610709b3
000822dc
07b46107
645460c7
74dc60e7
0df3000a
92dc6127
61470008
000a04dc
04c31173
0b58b2bc
1407045c
74dc0007
60260009
1e95345c
1e24345c
0a8b333c
0050533c
04c302d3
0b787ebc
1407045c
53dc0007
a0c70008
345c0c94
341c1e24
67f20400
76bc04c3
a0a60ba0
a02602d2
1e69345c
e87435e4
345c6046
345c1e95
341c1e44
60070004
40666c94
1e95245c
345c6086
345c1e95
341c1e24
68d20003
4cbc04c3
045c0b5b
00071407
40a65894
1e95245c
1e24345c
0400341c
04c368f2
0b6d66bc
1407045c
49940007
345c60c6
345c1e95
341c1e24
68d20003
e2bc04c3
045c0b7f
00071407
40e63a94
1e95245c
6abc04c3
045c0b5d
00071407
61063094
1e95345c
fcbc04c3
045c0b5c
00071407
41262694
1e95245c
04c30113
0b787ebc
1407045c
1b740007
1e69345c
f63560a7
345c6146
714c1e95
04c369d2
3664316c
04150007
1407045c
345c0153
341c1e24
67f24000
7cbc04c3
00730b68
00531fe6
01960026
08040c56
40c31016
1e24305c
0010341c
64f25fe6
0ba1a6bc
345c20c3
341c1e24
65d20010
d8bc04c3
20c30ba2
085602c3
00000804
1f36f016
70c3fc96
b2c351c3
000783c3
000bd2dc
a2dc2007
6007000b
000b72dc
0500a33c
133c0ac3
2ac3384e
0ac9dabc
000760c3
000ab4dc
10f8c01c
0000c11c
640c1cc3
04068c0c
44c616c3
69ac301c
0017311c
90c34664
82dc0007
bf5c0009
40260007
9f5c4077
c0f70047
101c08c3
111c68cc
2ac30017
b8bc35c3
50c30ba0
0dd40007
640c1cc3
09c38c4c
44c616c3
69ac301c
0017311c
0f134664
301c08c3
311c1498
2c0c0000
2abc40e6
01640892
3c0c0cf2
10fc301c
0000311c
5c4c6c0c
0007af5c
02d38ecc
301c08c3
311c149c
2c0c0000
2abc4186
01640892
3c0c0ff2
10fc301c
0000311c
5c4c6c0c
0007af5c
01c38eec
466439c3
08c350c3
1480301c
0000311c
41662c0c
08922abc
05f20164
5c4c7c0c
03d32206
301c08c3
311c1484
2c0c0000
2abc4166
01640892
7c0c05f2
23065c4c
08c301f3
1488301c
0000311c
41662c0c
08922abc
0df20164
5c4c7c0c
20372406
0027af5c
13c303c3
04bc39c3
50c30b26
10f8301c
0000311c
8c4c6c0c
200609c3
301c44c6
311c69ac
46640017
a5d20026
bf8705c3
1fe60254
f8760496
08040f56
3f36f016
00b7fa96
a2c32077
cf5c6037
40e70244
40e74054
a31c12d4
31540002
0002a31c
0ac305d4
17540007
a31c0b93
1d540003
0004a31c
01f35694
53544147
07d44147
31544107
0009a31c
06f34c94
3f544167
479441c7
1424301c
0000311c
301c0c10
311c1428
08d30000
143c301c
0000311c
301c0c10
311c1440
07930000
1434301c
0000311c
301c0c10
311c1438
06530000
142c301c
0000311c
301c0c10
311c1430
05130000
1464301c
0000311c
301c0c10
311c1468
03d30000
145c301c
0000311c
301c0c10
311c1460
02930000
146c301c
0000311c
301c0c10
311c1470
01530000
1444301c
0000311c
301c0c10
311c1448
2c100000
144c701c
0000711c
1454601c
0000611c
145c501c
0000511c
1458d01c
0000d11c
1450b01c
0000b11c
18c30097
b4bc4057
40c30892
32940007
0001a31c
201c2f94
211c1444
680c0000
80e403c3
1c100594
24101bc3
5c0cfd53
83e432c3
18100594
20100dc3
380cfc53
82e421c3
14100794
1460301c
0000311c
140c01f3
81e410c3
001724dc
1464201c
0000211c
301c0810
311c1468
2c100000
8007f913
001642dc
d0c30097
d0840057
0ebc08c3
03640892
703c1000
7de40010
001591dc
61476008
7c080754
0020703c
a4dc6147
a31c000a
0f940001
4dd244d7
301c4006
311c145c
0c0c0000
81e410c3
2ac30294
4c0f64d7
00e04f3c
101c04c3
111c68e4
41460017
08cbe6bc
14c307c3
b4bc4a06
40c30892
0007b0c3
101c6354
111c68d0
4a060017
0892b4bc
0df250c3
101c04c3
111c68d4
4a060017
0892b4bc
000750c3
001172dc
00070cc3
001132dc
101c05c3
111c68d8
4a060017
0892b4bc
000770c3
001072dc
41dc50e4
101c0010
111c68dc
4a060017
0892b4bc
9ea060c3
15c30cc3
b0bc24c3
600608cb
6a212cc3
05000c3c
0010173c
b0bc4406
caf208cb
101c07c3
111c68e0
4a060017
0892b4bc
c00760c3
000df2dc
c9dc67e4
373c000d
79a00010
678f1cc3
215c4026
005303c5
7808c025
fd5461a7
fb546147
b01c76c3
00970001
405719c3
0892b4bc
07f240c3
40072cc3
000bf2dc
03d36057
0ebc09c3
03640892
0de41000
20c31934
008f323c
03946147
025302c3
06342de4
61476808
00450394
2cc30173
42dc4007
303c000a
00970020
6baf6c20
1cc313b3
409724d2
67af6120
605793a0
40e403c3
000936dc
07dc8007
00170009
2ac314c3
24bc6457
50c30ba0
93dc0007
60170008
36c3cc0c
14c307c3
044f233c
0ac768bc
600730c3
301c7974
311c144c
2c0c0000
82e421c3
3bc30d94
180c6bf2
c4bc384c
50c30ab8
6b74a007
5bc3b84f
1bc30d13
301c29f2
311c1454
4c0c0000
80e402c3
1cc35d94
58542007
600767ec
6f8c5554
52546007
10f8901c
0000911c
680c29c3
0a068c0c
44c62457
69c8301c
0017311c
70c34664
0007b066
1cc34254
8f8c67ec
40062a06
46646fac
301c40c3
311c1454
4c0c0000
80e402c3
180c1794
27c3384c
f6bc34c3
50c30ac5
640c19c3
07c38c4c
44c62006
69c8301c
0017311c
a0074664
b84f1e74
06c30373
24c317c3
dcbc3cc3
50c30ba3
600c09c3
07c38c4c
44c62457
69c8301c
0017311c
a0274664
00d30894
fe8c501c
bf860093
a0060053
069605c3
0f56fc76
00000804
1478301c
0000311c
6ff26c0c
0b23bcbc
ff1c301c
21940007
147c001c
0000011c
0b23c6bc
18940007
147c001c
0000011c
0b23cabc
10940007
1478301c
0000311c
40254c0c
001c4c0f
011c147c
ccbc0000
60260b23
72c60053
080403c3
40c3f016
01c371c3
0ba070bc
14c350c3
19548007
0500643c
cabc06c3
20060b23
11940007
5a1d443c
07c30133
0340143c
eabc4286
03d208cb
98f2924c
ccbc06c3
14c30b23
0f5601c3
00000804
0136f016
81c360c3
70bc01c3
50c30ba0
0500763c
cabc07c3
80060b23
12940007
5a1d463c
08c30173
0340143c
eabc4286
03f208cb
00738026
96f2924c
ccbc07c3
04c30b23
0f568076
00000804
40c3f016
72c361c3
0ebc01c3
50c30892
04c35364
1554a007
780801d3
099432e4
16c304c3
eabc25c3
03f208cb
013304c3
ffe58025
041475e4
40075008
0006ef94
08040f56
40c33016
ff53001c
11548007
0500543c
cabc05c3
20c30b23
49f212c6
216604c3
0aa71cbc
ccbc05c3
00260b23
08040c56
50c33016
1d540007
04d201ac
b6bc2026
05c30b9f
556c2166
0aa71cbc
0500053c
0b23c8bc
10f8301c
0000311c
8c4c6c0c
356c05c3
301c4326
311c69dc
46640017
08040c56
50c33016
10f8301c
0000311c
8c0c6c0c
15c30c06
301c4326
311c69f4
46640017
000740c3
20061754
b0bc4c06
043c0891
c6bc0500
06d20b23
94bc04c3
80060ba7
301c0133
345c0080
638602e6
02f6345c
04c3b16f
08040c56
b6bc0006
08040ba7
60c37016
1e540007
a007a00c
746c1b54
05946027
344c140c
0b06b8bc
740f6006
301c744f
311c10f8
6c0c0000
05c38c4c
548c342c
6a10301c
0017311c
40064664
0e56580f
00000804
ff961016
001c40c3
8007ff53
345c2654
6dd20621
4741345c
69f26037
0e80043c
0ba7e6bc
00013f5c
0625345c
0629345c
043c68d2
e6bc0f00
60060ba7
062d345c
345c0026
69d20631
0ec0043c
0ba7e6bc
345c6006
00260635
08560196
00000804
0f36f016
80c3ff96
a2c3b1c3
241063c3
10f8301c
0000311c
8c0c6c0c
0408001c
44c62006
69d4301c
0017311c
50c34664
20373066
92dc0007
29c3000d
484c280c
716c48c3
0ab0fcbc
208605c3
38c326c3
0ac32ebc
c0070037
74ec1f54
0206331c
331c1054
18940285
235c38c3
400702e2
000b83dc
742c2364
30dc32e4
0193000b
235c38c3
400702f2
000a93dc
742c2364
40dc32e4
4017000a
74dc4007
255c0008
4f5c1819
34c30001
0001a31c
60260254
43f23264
76946007
09944027
155c68d2
31c31843
0004341c
6c546007
2d80753c
17c308c3
0ba734bc
67940007
096c28c3
0aa6c8bc
05f240c3
fed1401c
0b1334c3
202f34ec
406f540c
600f742c
208f37cc
40af57ac
1829355c
155c614d
216d1821
40cf556c
60ef758c
0340603c
17c306c3
b0bc4286
043c08cb
153c0200
42860340
08cbb0bc
ffff301c
0000311c
1839155c
355c23d2
708e1843
524f4006
57af540f
558f556f
70bc06c3
60c30ba0
0500783c
cabc07c3
00070b23
38c31594
6a1d333c
18c3724f
6b9d413c
ccbc07c3
28c30b23
60076a0c
49c31254
304c100c
36642ac3
04c30193
296c28c3
0aa6e8bc
603772c6
101c0093
2037fe9b
64bc05c3
301c0aa3
311c10f8
6c0c0000
05c38c4c
44c62006
69d4301c
0017311c
0bc34664
0ba7e6bc
4bf24017
60376026
101c0113
fc93fe66
fe67301c
fc336037
01960017
0f56f076
00000804
3f36f016
70c3e096
d2c32137
bf5c60f7
20060584
27b727f7
81d003d2
cbc300d3
43d22bc3
8d303bc3
22d22b57
40d7a411
7fe532c3
6047df66
003645dc
0b0d373c
133c7fe5
2177f88c
0b0d3b3c
133c7fe5
21b7f88c
46d24157
ff53601c
14dc2007
501c0035
511c10f8
740c0000
001c8c0c
1cc30080
301c44c6
311c699c
46640017
000780c3
0033b2dc
305c6006
e3ef03c5
23af2006
07c04f3c
32c340d7
44dc6027
cf5c0010
8f5c0007
3f3c0027
60b70780
1dc30117
34c34ad7
0ba4a6bc
2b5760c3
28c324d2
440f4bac
83dcc007
2b97000e
42dc2007
4ad70010
04dc4007
38c30010
9de42fb0
000fb8dc
09a40dc3
08d40027
21f72ad7
42374026
0240af3c
02370fd3
10f8501c
0000511c
8c0c740c
40861cc3
699c301c
0017311c
a0c34664
61f76026
6b940007
8c4c740c
1cc308c3
301c44c6
311c699c
46640017
07c00f3c
0ba7e6bc
20065bb3
28c32777
cf5c2baf
8f5c0007
3f3c0027
60b70780
01c32117
1dc30984
400619a4
07403f3c
0ba4a6bc
000760c3
67572794
74000c4c
21c32217
053532e4
601c8026
0393ff7c
2e803ac3
0b3ef4bc
0030453c
1ac36757
2c0c0600
b0bc4c4c
675708cb
b1004c4c
4fac38c3
80269284
26d22b57
640c2b57
640f6d00
0f3c8026
e6bc0740
631c0ba7
0394fe8c
1a948007
1615c007
200721d7
301c6154
311c10f8
6c0c0000
0ac38c4c
40861cc3
699c301c
0017311c
0a534664
45c3a006
9de4f473
a007a174
3bc33854
1f546007
0629135c
0b3c25d2
e6bc0f00
0b3c0ba7
15c30f00
3cc34006
0ba024bc
000760c3
2bc32594
0784325c
1ac30c0c
b0bc25c3
202608cb
135c3bc3
0313062d
1554e007
0280473c
e6bc04c3
04c30ba7
2bc315c3
24bc3cc3
60c30ba0
7d4c09f2
1ac30c0c
b0bc25c3
005308cb
41d7c006
301c4fd2
311c10f8
6c0c0000
0ac38c4c
40861cc3
699c301c
0017311c
c0074664
301c2115
311c10f8
6c0c0000
04c30b73
4ad71dc3
24bc3cc3
60c30ba0
0c150007
8c4c740c
1cc308c3
301c44c6
311c699c
46640017
67d74353
21170c0c
b0bc2dc3
28c308cb
03c1225c
4a544007
13c360d7
46542027
10f8301c
0000311c
8c0c6c0c
1cc30a06
301c44c6
311c699c
46640017
d06650c3
13540007
4ff24157
8dd29f8c
7fac2a06
30c34664
15c307d7
38c323c3
0ba3dcbc
007360c3
ff50601c
10f8901c
0000911c
640c19c3
05c38c4c
44c61cc3
699c301c
0017311c
c0274664
19c31154
8c4c640c
1cc308c3
301c44c6
311c699c
46640017
07c00f3c
0ba7e6bc
301c38d3
311c10f8
6c0c0000
08c38c4c
44c61cc3
699c301c
0017311c
4ad74664
608732c3
4f3c1794
215707c0
04c327d2
0ba7e6bc
ff53601c
1d8c3553
275c6157
42f201e9
14c36026
3abc4026
60c30ba8
6ad733d3
1c946007
20071bc3
215c1054
45d20621
0e800b3c
0ba7e6bc
3bc327d7
0747135c
235c4026
05d30625
2c54e007
0240073c
0ba7e6bc
7d2f67d7
2ad704b3
402721c3
3bc31b94
10546007
0631135c
0b3c25d2
e6bc0ec0
67d70ba7
325c2bc3
20260767
0635125c
eed201f3
02c0073c
0ba7e6bc
5d6f47d7
0f3c00f3
e6bc07c0
df060ba7
6ad72b93
202713c3
0009b4dc
32c340d7
62dc6067
a7970009
5194a007
301ca777
311c10f8
6c0c0000
001c8c0c
1cc30098
301c44c6
311c699c
46640017
000780c3
001392dc
f4bc15c3
60c30b1c
20940007
0c0c67d7
07401f3c
6c4c28c3
0abeb4bc
2ad705d2
56c327b7
08c30273
0b1c4cbc
46d22bc3
1ed2325c
077403e4
e7d20113
0282375c
031503e4
fe67601c
08c3a026
0b1ce6bc
10f8301c
0000311c
8c4c6c0c
1cc308c3
301c44c6
311c699c
46640017
34dcc007
a0070010
000ff4dc
67776006
02404f3c
6cbc04c3
67d70ace
1f3c0c0c
24c30740
a4bc6c4c
05d20ab1
b6bc04c3
0bb30ad2
29d21bc3
72bc04c3
20c30ace
315c1bc3
01131ee2
04c3efd2
0ace72bc
375c20c3
23e40292
04c30715
0ad2b6bc
fe66601c
0f3c1a53
b6bc0240
40260ad2
e4d247b7
375c6026
1bc30245
42dc2007
315c000c
7a721e24
1e27315c
4ad717b3
a4dc4007
801c000b
811c10f8
18c30000
8c0c640c
0408001c
44c61cc3
699c301c
0017311c
50c34664
42dc0007
67d7000a
4c4c2c0c
fcbc3cc3
05c30ab0
f4bc2ad7
00070abd
18c30e15
8c4c640c
1cc305c3
301c44c6
311c699c
46640017
11b3df86
321c74cc
60c7fdf8
202613b4
300d313c
0071341c
e4d26dd2
275c4026
3bc3023d
335c67d2
79721e24
315c1bc3
ebd21e27
19a4255c
74ec5f4f
0206331c
40260494
0225275c
6fd23bc3
19a4155c
1fe7135c
331c74ec
07940206
315c1bc3
75721e24
1e27315c
331c74ec
21540206
0285331c
41973e94
1bc34cf2
1e24315c
0040341c
015c66f2
00071ed2
05f30c15
2f54e007
01e9275c
2b944007
0282075c
25740007
236420c3
32e4742c
04332014
4cf24197
315c1bc3
341c1e24
66f20040
1ee2015c
0b150007
e00701f3
275c1254
4ff201e9
0292075c
06740007
236420c3
32e4742c
601c0634
0073fe66
fe67601c
64bc05c3
301c0aa3
311c10f8
6c0c0000
05c38c4c
44c61cc3
699c301c
0017311c
c4d24664
d0660093
c0260053
209606c3
0f56fc76
00000804
0736f016
90c3fb96
62c381c3
800673c3
54c304c3
0100af3c
40060373
63574137
43976037
af5c4077
60060047
09c360f7
2a0028c3
37c35a20
0ba934bc
03740007
0093a026
60076117
611705f4
46e49180
a2d2e574
05960026
0f56e076
00000804
fd963016
207740c3
53c302c3
1d548007
1b542007
19744007
60b76046
4000101c
0b9feebc
47a3145c
0b9feebc
3f3c20c3
60370080
1f3c04c3
35c30040
0b79febc
05150007
00731fe6
ff53001c
0c560396
00000804
eabc6006
08040bac
ff963016
000740c3
305c4154
341c1e44
60070002
105c3d94
21c31e24
8000501c
0005511c
40072583
20261594
0b59c0bc
1407045c
2a740007
1e24345c
345c7272
a0061e27
0002511c
00463583
21546007
400603f3
0006211c
a0061283
0004511c
12e425c3
1f3c1394
23c30030
0bad14bc
0c740007
1e24345c
511ca006
35830002
40a668d2
1407245c
1fe60073
00260053
0c560196
00000804
0ad21016
400729d2
babc0774
00070b5a
1fe60515
001c0073
0856ff53
00000804
600c05d2
5cbc2dcc
08040b84
50c33016
2d540007
6ed26029
03d2002c
0bad74bc
08d2148c
1118301c
0000311c
6e0c6c0c
144c3664
301c0ed2
311c10f8
6c0c0000
20068c4c
301c4286
311c6988
46640017
10f8301c
0000311c
8c4c6c0c
200605c3
301c4286
311c6988
46640017
0c560006
00000804
50c33016
000740c3
301c1c54
311c10f8
6c0c0000
001c8c0c
35cc0920
301c4226
311c6a24
46640017
0bd240c3
b2bc15c3
00070b6b
04c30615
5cbc35cc
80060b84
0c5604c3
00000804
0136f016
601c70c3
0007ff53
801c2654
811c10f8
28c30000
8c0c680c
3dcc0206
301c4406
311c6a30
46640017
d06650c3
13540007
0b1c16bc
0dd260c3
680c28c3
05c38c4c
44063dcc
6a30301c
0017311c
00734664
c026bc2f
807606c3
08040f56
2cbc03d2
08040b84
0136f016
71c360c3
1478301c
0000311c
adf2ac0c
0ba6e0bc
09540027
3154c007
10f8301c
0000311c
04336c0c
2954c007
10f8801c
0000811c
680c28c3
001c8c0c
17c30098
301c4246
311c6a44
46640017
0bd250c3
27c316c3
0b8476bc
12150007
02bc05c3
01b30bae
680c28c3
06c38c4c
416617c3
6a44301c
0017311c
00534664
05c3a006
0f568076
00000804
06bc2006
08040bae
ff96f016
51c340c3
73c362c3
0a759abc
3f5c0037
69d20001
15c304c3
37c326c3
0afbd4bc
02f27fe6
03c36006
0f560196
00000804
0af574bc
1fe630c3
03c362f2
00000804
0aefaabc
1fe630c3
03c362f2
00000804
0ae698bc
1fe630c3
03c362f2
00000804
0ae67abc
1fe630c3
03c362f2
00000804
0ae55abc
00000804
0ae542bc
00000804
0ae4e8bc
1fe630c3
03c362f2
00000804
0ae318bc
00000804
60c3f016
42c371c3
0ae318bc
88d250c3
32c3500c
043503e4
1fe6100f
06c30193
60bc17c3
30c30af2
65f21fe6
83d204c3
03c3b00f
08040f56
40c31016
7ebc0cd2
301c0ae2
311c1110
6c0c0000
07c4335c
366404c3
08040856
501c3016
511c1110
740c0000
0784335c
36640206
0ad240c3
0ae25ebc
740c07d2
07c4335c
366404c3
04c38006
08040c56
00180005
73206f6e
6f707075
66207472
6520726f
726f7272
72747320
73676e69
69756220
6920746c
0000006e
43414843
00004148
00004345
004d4343
004c4c41
0000003a
00485351
53444345
00000041
00484441
004b5350
2d344352
00414853
2d344352
0035444d
2d534544
33434243
4148532d
00000000
31534541
532d3832
00004148
32534541
532d3635
00004148
2d454844
2d415352
31534541
532d3832
00004148
2d454844
2d415352
32534541
532d3635
00004148
31534541
432d3832
382d4d43
00000000
32534541
432d3635
382d4d43
00000000
48444345
43452d45
2d415344
31534541
432d3832
00004d43
48444345
43452d45
2d415344
31534541
432d3832
382d4d43
00000000
48444345
43452d45
2d415344
32534541
432d3635
382d4d43
00000000
48444345
53522d45
45412d41
38323153
4148532d
00000000
48444345
53522d45
45412d41
36353253
4148532d
00000000
48444345
43452d45
2d415344
31534541
532d3832
00004148
48444345
43452d45
2d415344
32534541
532d3635
00004148
48444345
53522d45
43522d41
48532d34
00000041
48444345
53522d45
45442d41
42432d53
532d3343
00004148
48444345
43452d45
2d415344
2d344352
00414853
48444345
43452d45
2d415344
2d534544
33434243
4148532d
00000000
31534541
532d3832
35324148
00000036
32534541
532d3635
35324148
00000036
2d454844
2d415352
31534541
532d3832
35324148
00000036
2d454844
2d415352
32534541
532d3635
35324148
00000036
48444345
4153522d
5345412d
2d383231
00414853
48444345
4153522d
5345412d
2d363532
00414853
48444345
4443452d
412d4153
32315345
48532d38
00000041
48444345
4443452d
412d4153
35325345
48532d36
00000041
48444345
4153522d
3443522d
4148532d
00000000
48444345
4153522d
5345442d
4342432d
48532d33
00000041
48444345
4443452d
522d4153
532d3443
00004148
48444345
4443452d
442d4153
432d5345
2d334342
00414853
31534541
472d3832
532d4d43
35324148
00000036
32534541
472d3635
532d4d43
38334148
00000034
2d454844
2d415352
31534541
472d3832
532d4d43
35324148
00000036
2d454844
2d415352
32534541
472d3635
532d4d43
38334148
00000034
48444345
53522d45
45412d41
38323153
4d43472d
4148532d
00363532
48444345
53522d45
45412d41
36353253
4d43472d
4148532d
00343833
48444345
43452d45
2d415344
31534541
472d3832
532d4d43
35324148
00000036
48444345
43452d45
2d415344
32534541
472d3635
532d4d43
38334148
00000034
48444345
4153522d
5345412d
2d383231
2d4d4347
32414853
00003635
48444345
4153522d
5345412d
2d363532
2d4d4347
33414853
00003438
48444345
4443452d
412d4153
32315345
43472d38
48532d4d
36353241
00000000
48444345
4443452d
412d4153
35325345
43472d36
48532d4d
34383341
00000000
48444345
53522d45
45412d41
38323153
4148532d
00363532
48444345
43452d45
2d415344
31534541
532d3832
35324148
00000036
48444345
4153522d
5345412d
2d383231
32414853
00003635
48444345
4443452d
412d4153
32315345
48532d38
36353241
00000000
48444345
53522d45
45412d41
36353253
4148532d
00343833
48444345
43452d45
2d415344
32534541
532d3635
38334148
00000034
48444345
4153522d
5345412d
2d363532
33414853
00003438
48444345
4443452d
412d4153
35325345
48532d36
34383341
00000000
2d484441
31534541
532d3832
00004148
2d484445
2d415352
2d534544
33434243
4148532d
00000000
646e6553
76726553
654b7265
63784579
676e6168
00000065
65657246
4579654b
61686378
0065676e
646e6553
74726543
63696669
56657461
66697265
00000079
36363636
36363636
36363636
36363636
36363636
36363636
36363636
36363636
36363636
36363636
36363636
36363636
5c5c5c5c
5c5c5c5c
5c5c5c5c
5c5c5c5c
5c5c5c5c
5c5c5c5c
5c5c5c5c
5c5c5c5c
5c5c5c5c
5c5c5c5c
5c5c5c5c
5c5c5c5c
6c697542
35444d64
7265435f
72655674
00796669
6c697542
41485364
7265435f
72655674
00796669
646e6553
65696c43
654b746e
63784579
676e6168
00000065
646e6553
65696c43
6548746e
006f6c6c
00175e1c
00175e24
00175e2c
00175e3c
00175e48
00175e54
00175e68
00175e7c
00175e8c
00175e9c
00175eb4
00175ed0
00175eec
00175f04
00175f1c
00175f34
00175f4c
00175f60
00175f78
00175f8c
00175fa8
00175fb8
00175fc8
00175fe0
00175ff8
0017600c
00176020
00176038
00176050
00176064
0017607c
00176090
001760a8
001760bc
001760d0
001760ec
00176108
00176124
00176140
00176160
00176180
0017619c
001761b8
001761d8
001761f8
00176210
0017622c
00176244
00176260
00176278
00176294
001762ac
001762c8
001762d8
00000005
00000004
0000000a
0000002f
00000035
00000033
00000039
000000a0
000000a1
000000ac
000000ae
000000af
00000013
00000014
00000009
0000000a
00000011
00000012
00000007
00000008
0000003c
0000003d
00000067
0000006b
0000000e
0000000f
00000004
00000005
0000000c
0000000d
00000002
00000003
0000009c
0000009d
0000009e
0000009f
0000002f
00000030
0000002b
0000002c
00000031
00000032
0000002d
0000002e
00000027
00000023
00000029
00000025
00000028
00000024
0000002a
00000026
00000034
00000016
646e6553
74726543
63696669
00657461
544e4c43
52565253
6c697542
6e694664
65687369
00000064
6c697542
35444d64
00000000
6c697542
41485364
00000000
61486f44
6853646e
4d656b61
00006773
65536f44
72657672
4579654b
61686378
0065676e
65536f44
6f697373
6369546e
0074656b
65436f44
66697472
74616369
00000065
6c436f44
746e6569
4579654b
61686378
0065676e
65436f44
66697472
74616369
72655665
00796669
79706f43
6f636544
54646564
3035586f
00000039
776f7247
7074754f
75427475
72656666
00000000
776f7247
75706e49
66754274
00726566
69726853
6e496b6e
42747570
65666675
00000072
69726853
754f6b6e
74757074
66667542
00007265
65657246
004c5353
65657246
646e6148
6b616873
73655265
6372756f
00007365
5f4c5353
6f736552
65637275
65657246
00000000
65657246
61727241
00007379
74696e49
004c5353
65657246
39303558
00000000
65657246
39303558
656d614e
00000000
65657246
68706943
00737265
65657246
5f4c5353
00787443
5f4c5353
52787443
756f7365
46656372
00656572
00000041
00004242
00434343
44444444
00000000
45454545
00000045
46464646
00004646
47474747
00474747
48484848
48484848
00000000
49494949
49494949
00000049
656b614d
4d6c7353
65747361
63655372
00746572
69726544
654b6576
00007379
4b746553
00737965
58534c54
6572465f
6c6c4165
00000000
58534c54
77654e5f
00000000
58534c54
7365535f
6e6f6973
6b636954
465f7465
00656572
58534c54
7365535f
6e6f6973
6b636954
435f7465
74616572
00000065
58534c54
6573555f
4678614d
6d676172
00746e65
7473616d
73207265
65726365
00000074
69726544
6c546576
79654b73
00000073
2079656b
61707865
6f69736e
0000006e
544e4c43
65696c63
6620746e
73696e69
00646568
76726573
66207265
73696e69
00646568
00465250
61685f70
00006873
52506f64
00000046
63656843
73634f6b
71655270
74736575
00000000
4f746547
45707363
7972746e
00000000
4f746547
53707363
75746174
00000073
63656843
7265436b
53434f74
00000050
65657246
5053434f
00000000
65657246
7073634f
72746e45
00000079
454e4f4e
00000000
0035444d
00534544
00534541
0000002c
0000000d
0000000a
636f7250
7079542d
00000065
2d534541
2d383231
00434243
2d534541
2d323931
00434243
2d534541
2d363532
00434243
2d534541
2d383231
00525443
2d534541
2d323931
00525443
2d534541
2d363532
00525443
2d534544
00434243
2d534544
33454445
4342432d
00000000
0000000b
00000007
0000000c
65747845
6c616e72
65657246
39303558
00000000
666c6f77
5f4c5353
5f505645
65747942
4b6f5473
00007965
666c6f77
5f4c5353
5f4f4942
65657266
00000000
636f7250
42737365
65666675
00000072
666c6f77
5f6c7373
72636564
5f747079
66667562
6b5f7265
00007965
546d6550
7265446f
00000000
43646441
00000041
666c6f77
5f4c5353
74726543
616e614d
46726567
00656572
666c6f77
5f4c5353
74726543
616e614d
4e726567
655f7765
00000078
65657246
00726544
6f6c6c41
72654463
00000000
666c6f77
5f4c5353
0077656e
666c6f77
5f4c5353
5f585443
5f77656e
00676e72
666c6f77
5f4c5353
5f585443
5f77656e
00007865
000620c3
31c32829
31a32849
31a32809
31a32869
31a32889
31a328a9
002662f2
00000804
0804002c
0804004c
40a1041c
002602d2
00000804
0542041c
002602d2
00000804
40c31016
0bb542bc
07f26026
48bc04c3
02d20bb5
30c30026
085603c3
00000804
40c31016
0bb54ebc
03f26026
090b343c
085603c3
00000804
305c20c3
6c6c0744
63d21fe6
36640bac
00000804
305c20c3
6dec0744
63d21fe6
36640bac
00000804
00000804
08040006
08040006
08040006
632cff96
03546087
03946207
02530006
0f946107
0dd2026c
63ec4006
0003341c
402662f2
0016123c
0f5c2037
00530001
01960026
00000804
08040006
205c6006
43d20ca4
00d30026
00856025
f8946087
080402c3
60c37016
315c41c3
60070d64
674c2394
0200341c
1e946007
a4bc01c3
02d20bb5
50c30026
303c134c
66d20084
341c73ec
62d20003
4ebca026
02d20bb5
365ca026
03c302b3
0010041c
a2f206f2
50c30026
a0260053
0e5605c3
00000804
05f220c3
408500f3
045401e4
1cf2080c
00260053
00000804
09b3031c
021c09d4
20a6f694
0a7c5cbc
0010303c
600600d3
09b4031c
61c60294
080403c3
61ac20c3
0001341c
67d20026
6ac90006
00ff331c
00260294
00000804
40c33016
12c301c3
a1224006
b12235c3
a5223503
63d23583
00b30006
40c74025
0026f594
08040c56
70c3f016
41c362c3
0193a006
17c304c3
0060243c
0bb60abc
03d28185
00b30026
56e4a025
0006f414
08040f56
00870364
00c70354
00260394
303c00d3
7fe50076
f88c033c
00000804
00000804
00000804
00000804
70c3f016
301c61c3
311c10fc
6c0c0000
30c98c0c
30e921c3
412c313c
323c5109
312981ac
c1ac313c
0bb460e7
345c6006
043c07cd
20060fa0
a4bc40c6
03930bce
0200563c
143c05c3
40c60300
0bcdd2bc
14540007
063c7e6c
2c8c02c0
d2bc4cac
0cf20bcd
145c2026
043c07cd
15c30fa0
b4bc40c6
00260bcd
00060053
08040f56
1f36f016
91c380c3
e44c842c
54c30653
009e253c
0020623c
2ed467e4
331c7009
0d9400dd
0b3540a7
0020043c
f7c4101c
0017111c
d2bc40c6
07d20bcd
66077009
74091694
13356027
111c501c
0000511c
6dac740c
015c18c3
14c30784
366426c3
740c0bf2
08c36d8c
02b33664
9300ff20
e02783d2
59c3cdd4
6dd2742c
111c301c
0000311c
6dac6c0c
015c18c3
20060784
366421c3
111c401c
0000411c
335c700c
28c30da4
0784025c
346c59c3
3664548c
19c3b4ac
c00664d0
c4c3a6c3
45c30753
009e243c
0020723c
37d47be4
20071ac3
74091c94
00dd331c
40a71894
053c1635
101c0020
111cf7c4
40c60017
0bcdd2bc
1cc30cf2
6dcc640c
025c28c3
15c30784
366427c3
0001a01c
1194c007
66077409
70090e94
0b356027
640c1cc3
28c36dec
0784025c
27c315c3
c0263664
b780b7a4
b31ca4d2
c4d40001
a0075ac3
19c31094
6dd264ac
111c301c
0000311c
6dcc6c0c
025c28c3
1ac30784
36642ac3
1094c007
74ac59c3
301c6dd2
311c111c
6c0c0000
18c36dec
0784015c
26c316c3
3ac33664
64d236a3
38c3a026
18c3aeaf
49d246cc
74ec59c3
23e466d2
08c30454
0bc14ebc
68ec29c3
6acf28c3
f8760006
08040f56
9ebc03ac
08040bc3
60c37016
0253a006
433c6c2c
01935a1d
14c306c3
0bd528bc
345c06f2
7fe50de4
0a356027
95f2902c
796ca025
12c34c4c
eb7451e4
04c38006
08040e56
fe963016
41c350c3
14542007
10a4315c
10546007
92bc0fc3
345c0bcd
001710a4
03f430e4
00f30c20
14c305c3
60bc4006
00060bd5
0c560296
00000804
40c33016
426c51c3
65d268ac
a6bc488c
0af20bcb
111c301c
0000311c
6d4c6c0c
15c304c3
0c563664
00000804
40c33016
0380503c
a0bc15c3
09f20bb7
4ebc04c3
04c30bc1
a0bc15c3
02d20bb7
0c56128f
00000804
e2967016
616c50c3
60276cac
626c1e94
1b546007
0bb7b6bc
6cac766c
70546007
05404f3c
14c305c3
0bb56abc
000720c3
766c6774
10c30cac
079421e4
2c8c04c3
0bcdd2bc
5c540007
ecbc05c3
60c30bd5
58540007
16c305c3
0bd528bc
52940007
153c05c3
90bc0380
00070bd5
05c34b94
58ac388c
0bd56abc
000740c3
05c34394
82bc16c3
00070bb7
1b4c3dd4
0bb55ebc
6a060ed2
3f3c6777
60370740
14c305c3
3f3c26c3
5ebc0040
01530bd6
111c301c
0000311c
6d0c6c0c
16c305c3
766c3664
36e46cd2
301c0a54
311c111c
6c0c0000
055c6d2c
366407a4
d66f966c
b6bc05c3
05c30bb7
6cbc366c
05c30be6
0bd858bc
21c3366c
045442e4
9abc05c3
00060be7
1fe60053
0e561e96
00000804
0136f016
60c3f096
005c41c3
805c0784
265c0c81
40071244
20071754
001822dc
111c301c
0000311c
68ac2c0c
510c6c0c
d04cb02c
0037100c
03c3860c
25c312c3
466436c3
301c2dd3
311c111c
6c0c0000
0dc4335c
70c33664
06c388d2
88bc14c3
00070bb6
0015e3dc
03a05f3c
15c306c3
0bb760bc
2d740007
20c606c3
0bd804bc
0380463c
14c305c3
d2bc40c6
00070bcd
04c35054
40c615c3
0bcdb4bc
03e0063c
40c62006
0bcea4bc
9cbc06c3
06c30be7
0bb586bc
e7f208d2
65f238c3
15c306c3
0bd470bc
cabc06c3
30c30bb7
0b156007
111c301c
0000311c
6e2c6c0c
206606c3
23f33664
60077a6c
4f3c1154
06c303a0
a0bc14c3
09f20bb7
4ebc06c3
06c30bc1
a0bc14c3
02d20bb7
796c1a8f
60276cac
365c1094
40060a04
0004211c
69d23283
111c301c
0000311c
6e4c6c0c
366406c3
0784065c
03a01f3c
0bf062bc
03d2186c
0bfafabc
fff0383c
f88c533c
0b0d373c
7f327fe5
438345c3
065c8bd2
200607a4
0bfab8bc
07a4065c
b2bc2006
1b2c0bfa
0bb548bc
e6d202f2
07a4065c
a2bc2006
065c0bfa
202607a4
0bfab8bc
365c6006
7b2c0867
09546087
07546207
6dd27a6c
0de4335c
09946027
c0bc06c3
06c30bd8
04bc2126
00f30bd8
06c386d2
40062146
0bd8d4bc
111c301c
0000311c
6e6c6c0c
366406c3
0a04365c
0084433c
1b2c85d2
0bb548bc
38c304f2
10546007
c0bc06c3
06c30bd8
04bc2126
065c0bd8
202607a4
0bfab2bc
2054a007
8bd20353
42bc1b2c
07d20bb5
07a4065c
b2bc2026
02930bfa
1254e007
c0bc06c3
06c30bd8
04bc2126
065c0bd8
202607a4
0bfab2bc
07a4065c
a2bc2026
365c0bfa
70920c84
0c87365c
0c04365c
3e546007
03000f3c
0bcd92bc
065c6317
4c200c24
165c6357
6ca00c44
07156007
101c5fe5
111c4240
6c80000f
21944007
869f201c
0001211c
30e402c3
763c1ad4
07c318c0
03a01f3c
d2bc40c6
00070bcd
465c1094
04c30c04
0bb540bc
04c350c3
0bb53ebc
06c330c3
25c317c3
0bd8fabc
0c04065c
0bcf06bc
165c2006
7b2c0c07
03546087
11946107
6fd27a6c
1f3c06c3
74bc0040
09f20bb5
00813f5c
65d26732
3a6c06c3
0bd414bc
1f3c06c3
1cbc03a0
18c30bc6
301c2cd2
311c111c
6c0c0000
065c6eac
163c0784
36644740
80761096
08040f56
40c3f016
72c361c3
0bc1dabc
0cf250c3
204604c3
0bd804bc
1f24345c
081b353c
1f27345c
602601d3
09e7345c
111c301c
0000311c
6d6c6c0c
16c304c3
366427c3
08040f56
0736f016
91c3fe96
1f5c2026
46460035
003d2f5c
0e9039c3
200718c3
305c5d54
600722a4
a05c5954
13c322c3
54c38006
323c0293
044c200c
6c2c6c00
069438e4
700c89d2
06946027
40250093
f27426e4
a02574c3
47c32705
05155ae4
c42c71c3
feb34006
3a548007
00607f3c
3c0909c3
0bc824bc
000760c3
20292954
821c81c3
a0460001
5aa20433
241c4037
023c007f
3f5c0057
30640001
15156007
04544fe7
4006306c
04c30193
0bb5fcbc
02d30cf2
333c708c
30e42a1d
40250654
f97421e4
0c5421e4
85e4a025
e025df15
00801f3c
72e421c3
0026cc94
00060053
e0760296
08040f56
0336f016
70c3f796
62c341c3
0bc788bc
48dc0007
b34c000b
4ebc05c3
801c0bb5
0ef20000
0044353c
345c69d2
6ca50d24
3a1d343c
0001801c
853c63f2
06c308cb
24bc2606
90c30bc8
341c738c
62d20002
e00603f2
29c308d3
13c36829
2f3c2045
c2bc0040
00070be0
18c33b94
60d727d2
0006341c
14dc6007
738c0008
32834057
2e546007
2097730c
60073183
732c2954
328340d7
24546007
2117734c
60073183
61571f54
0804133c
20072037
345c6694
60670e84
3f5c0d94
23c30001
335c7d6c
60470ea4
40260294
326432c3
361c00f3
333c0002
7fe50b0d
60077f32
e0264e54
101c06c3
111cf201
3cbc0050
60c30bc8
341c738c
60070001
00072554
e0252354
12c34029
2f3c2045
c2bc0040
00070be0
38c31994
60d766d2
0006341c
2d946007
2057738c
6ed23183
4097730c
6ad23283
20d7732c
66d23183
4117734c
60073283
b34c1c94
0084353c
c4f265d2
600739c3
738c1454
0003341c
05c367d2
0bb54ebc
07c303d2
05c3ebd2
0bb54ebc
0b0d303c
033c7fe5
0053f88c
09960026
0f56c076
00000804
3f36f016
70c3ff96
c3c352c3
20372a8c
101c02c3
111cf201
3cbc0050
b0c30bc8
b05c03d2
05c30009
24bc2606
40c30bc8
802902d2
101c05c3
111c9a12
3cbc506f
60c30bc8
c02602d2
0200853c
18c307c3
0bd32abc
0007a0c3
07c31054
0bc1dabc
0016303c
0b0d333c
233c33c4
1ac3f88c
32e4646c
000e36dc
6007766c
000df2dc
10fc301c
0000311c
2c0c6c0c
3051215c
341c32c3
6ad20010
121c08c3
40c60604
0bcdd2bc
a4dc0007
07c3000c
90bc18c3
00070bd5
000c34dc
02c0d53c
1dc307c3
6abc566c
00070bd5
000b94dc
34c390c3
32643ba3
901c63d2
4cc30001
b9a3b6c3
c0261533
25f219c3
62d270ac
63c36026
14c307c3
0bd528bc
b4dc0007
07c30009
82bc14c3
00070bb7
000946dc
eabc0017
09d20bb5
0650303c
7d806212
60276c28
000882dc
233c734c
46d20a4b
64d23ac3
60076c6c
39c37ed4
70ac6fd2
17946007
14c307c3
3ebc25c3
303c0bc7
7fe50b0d
63837f52
4bd20193
68f270ac
14c307c3
3ebc25c3
69c30bc7
c02602f2
6ad2718c
68f270ac
143c08c3
40c60180
0bcdd2bc
ccd20dd2
30ac566c
23e431c3
0dc35294
d2bc308c
00070bcd
718c4c94
08c369d2
0180143c
d2bc40c6
00070bcd
512c4294
08c347d2
1ebc310c
00070bb6
516c3a94
08c347d2
1ebc314c
00070bb6
07c33254
25c314c3
0bba78bc
2b540007
27f21bc3
341c734c
6007020c
01932454
4ad229c3
4ebc134c
06f20bb5
a4bc04c3
00070bb5
05c31894
b0bc14c3
00070bb5
155c1254
31c302b3
0002341c
045c6cf2
368c0f64
0bb5debc
07c306d2
06bc15c3
07f20bba
8007902c
fff574dc
80060053
019604c3
0f56fc76
00000804
3f36f016
50c3fb96
c2c3d1c3
10fc301c
0000311c
ec0c6c0c
075c0a06
355c09fd
c00607e4
612786c3
853c6294
46c30380
643c0853
355c100c
333c0684
033c4a1d
18c30200
d2bc40c6
00370bcd
32940007
0684355c
6f0c6f01
007703c4
1f5c178f
175c0021
2f5c0a15
275c0001
301c0a05
311c111c
4c0c0000
0684355c
4a8c6f01
0283035c
03642664
0a0d075c
1430073c
40c618c3
0bcdb4bc
0684355c
0e8c6f01
0bb5eabc
0650303c
75806212
14c3cc29
80250133
06a4355c
40e403c3
c006bb14
556c16c3
801c778c
425c0001
04c304a4
0d1530e4
0684355c
1a1d233c
1cc3766c
766c640f
123c05c3
0cd30530
09938006
100cb43c
0684355c
4a1d933c
431009c3
14c305c3
3dc329c3
0bbb3abc
040f1cc3
39540007
23c33ac4
08c36137
ccf20dd2
4d20778c
135c756c
01c30484
2b7420e4
175c2c06
2f5c09fd
275c0081
60060a15
0a05375c
111c401c
0000411c
355c500c
0bc30684
4a8c6c01
0283035c
03642664
0a0d075c
0684355c
6c811bc3
1430073c
0200133c
b4bc40c6
700c0bcd
00466ecc
03f33664
255c8025
32c306a4
b11443e4
48c398c3
15548007
111c301c
0000311c
6ecc6c0c
36640046
0cc3366c
766c200f
153c05c3
4c8c0380
a6bc6cac
90c30bcb
059609c3
0f56fc76
00000804
40c37016
305c61c3
60070684
305c2454
600706a4
03f31e94
04c36c2c
5a1d133c
5ebc26c3
00070bbc
a0251794
2c4c716c
52e421c3
345cf274
6dd20904
6bf2718c
debc04c3
345c0bd2
60250be4
0be7345c
fdb3a006
0e560006
00000804
70c3f016
0784005c
0be7e8bc
1b740007
453c57c3
02b35a4e
200604c3
0bc824bc
0ed260c3
260604c3
0bc824bc
08d230c3
0784075c
0200143c
c0bc26c3
900c0be8
eb9445e4
08040f56
0136f016
50c3ff96
62c381c3
0bc6dcbc
23540007
1884355c
05546067
19c4355c
11546007
111c301c
0000311c
335c6c0c
40060c24
02c34037
23c312c3
3cbc35c3
01330be5
111c301c
0000311c
6eec6c0c
366405c3
07931fe6
6007762c
783c2594
07c30200
0380153c
d2bc40c6
00070bcd
355c2e54
7f8507e4
16b46027
03e0453c
2cbc04c3
07f20bb5
14c307c3
d2bc40c6
0af20bcd
2cbc04c3
00070bb5
766c1854
62e423c3
05c31454
a2bc16c3
40c30bb5
05c307d2
40062146
0bb9e4bc
05c30113
26c318c3
0bd9f0bc
005304c3
01960006
0f568076
00000804
fd96f016
3f3c50c3
200600c0
fe7e133c
10fc201c
0000211c
880c480c
44bc13c3
00770bbd
3d540007
205705c3
48bc4097
40c30bb6
05c305f2
0bbd72bc
609723d3
12c3566c
135431e4
07e4355c
0f356067
2384355c
355c7972
301c2387
311c111c
6c0c0000
05c36e2c
36642066
205705c3
96bc4097
00070bbd
301c0f15
311c1110
6c0c0000
0684435c
20060286
60064b06
1fe64664
05c31eb3
0bbd72bc
1e130026
12c350c9
323c50e9
310940ac
81ac313c
323c5129
60e7c1ac
4a060535
09fd245c
6e6603d3
09fd345c
145c2c86
2f5c0a15
245c0021
345c0a0d
60370a01
0030341c
2f5c65d2
245c0001
60660a4d
0a05345c
1430043c
40c62006
0891b0bc
111c301c
0000311c
6ecc6c0c
36640046
0a01345c
06946067
0a49245c
09fd245c
60060093
09fd345c
145c2c86
40060a15
0a0d245c
0bc254bc
00070164
301c4854
311c111c
6c0c0000
36646f0c
3f940007
0bc27abc
00070164
30c93a94
30e921c3
412c313c
323c5109
312981ac
c1ac313c
063560e7
07c1345c
32dc6027
52660008
09fd245c
345c6066
2c860a05
0a15145c
245c4006
043c0a0d
20061430
a4bc40c6
301c0bce
311c111c
6c0c0000
00666ecc
301c3664
311c1110
6c0c0000
0684435c
20060286
60064326
0b734664
64bc05c3
20c30bb7
09d200b7
200605c3
0bd9f0bc
72bc05c3
09b30bbd
09a4655c
21c331c9
313c31e9
6027412c
145c1294
21c309b9
09c1145c
412c313c
09c9245c
81ac323c
09d1145c
c1ac013c
60c302d2
111c701c
0000711c
6f2c7c0c
366405c3
29540027
19c4355c
200605c3
d090201c
0003211c
10946007
2144355c
06d46007
debc05c3
40c30bc5
05c30ad2
201c2006
211ca120
e4bc0007
01b30bb9
6f4c7c0c
366405c3
05c308d2
24c316c3
0bb9e4bc
005304c3
03960006
08040f56
0136f016
81c340c3
1244705c
aabc2006
500c0bc1
0464125c
0014313c
2e546007
60076bcc
6aac2b94
28546007
1f24345c
0001341c
22946007
0584545c
1e94a007
353c31c3
325c081b
601c0467
611c111c
780c0000
6f6c500c
36640aac
0e940027
1f24345c
081b303c
1f27345c
6d6c780c
20a604c3
366425c3
345c0353
60921f24
1f27345c
e2d257c3
04c3a026
402618c3
0bc0d8bc
0df260c3
6cac716c
07546047
04c3a6f2
25c32026
0bb9e4bc
0e731fe6
10fc301c
0000311c
6c0c6c0c
21c32e49
313c2e69
6027412c
345c0f94
6cd20584
145c2006
04c30587
366416c3
40bc06c3
1fc60bd3
a9d20b13
1244045c
2384305c
1e546007
03933664
b8bc04c3
04c30be7
a2bc2026
04c30be7
0bb580bc
27d40007
6cac716c
06946047
debc04c3
00070bc5
04c31e54
84bc16c3
50c30bb5
06c306d2
0bd340bc
05f30006
66d2724c
15c304c3
0bd804bc
04c30193
0bd51cbc
0cf250c3
16c304c3
0bb582bc
06940027
40bc06c3
05c30bd3
301c0313
311c10fc
6c0c0000
2e496c0c
2e6921c3
412c313c
05946027
16c304c3
0bc690bc
40bc06c3
04c30bd3
0bbe02bc
0f568076
00000804
60c3f016
44bc71c3
00070bbf
365c2894
335c0744
60070a84
1bac2254
50c33664
1d540007
60076009
780c1a54
02b38c0c
125446e4
0744345c
0a84335c
13ac6dd2
10c33664
05c309d2
0bce28bc
04c305f2
44bc17c3
904c0bbf
eb948007
08040f56
0804002c
305c20c3
335c0744
1fe60dc4
0bac63d2
08043664
0bc044bc
1fe602d2
00000804
30c37016
0b8551c3
81004d2c
20290373
0020313c
19d432e4
331c6009
0f9400dd
0d352067
70126069
363cc049
40a9c1ac
c08932a3
41ac363c
085453e4
0020313c
50200180
e4d44027
0e560006
00000804
400c640c
28ec6cec
08040ca0
00000804
7cbc03ac
08040bc4
50c37016
63ec61c3
6cf28006
343c0253
57ec0067
16c30d00
d2bc40c6
09d20bcd
355c8025
23c30404
f21442e4
00530006
0e560026
00000804
0336f016
61c380c3
600763ec
80062a54
901c54c3
911c1110
03b30000
333c780c
08c34a1d
0530133c
0bc088bc
580c70c3
123c07d2
123c4a1d
a0255b9d
19c30173
335c640c
023c07c4
36644a1d
733c780c
80254b9d
43e4782c
35e4e214
b82f0254
0f56c076
00000804
0736f016
91c360c3
84bca2c3
50c30bc0
69540007
15c306c3
0bc0a4bc
debc06c3
06f20bc5
80f8701c
0017711c
301c00f3
311c111c
6c0c0000
140cec8c
301c0cd2
311c1110
6c0c0000
0864435c
4086342c
466437c3
1abc06c3
80060bc8
10fc801c
0000811c
1110701c
0000711c
740c0473
133c06c3
febc4a1d
18c30bcc
6c0c640c
12c34e49
323c4e69
602740ac
740c1254
133c06c3
2cbc4a1d
7c0c0bc6
335c540c
023c07c4
36644a1d
4006740c
4b9d233c
742c8025
41e413c3
06c3db14
2ac319c3
0bcc1cbc
10fc301c
0000311c
6c0c6c0c
12c34e49
323c4e69
602740ac
06c30454
0bc5eebc
e07605c3
08040f56
21c32006
0bc0d8bc
04d27fe6
0bd340bc
03c36006
00000804
41c33016
28d252c3
22bc12c3
14c30bcf
b4bc25c3
0c560bcd
00000804
0136f016
81c350c3
40bc012c
60c30bcf
35540007
05c0453c
f000152c
54c30493
009e253c
0020323c
20d431e4
331c7009
159400dd
13354067
70127069
303c1049
30a9c1ac
108931a3
41ac303c
079483e4
143c06c3
5f850060
0bc15abc
32c35409
91806045
20273e20
06c3dbd4
0bc042bc
05f240c3
06bc06c3
64c30bcf
807606c3
08040f56
305c1016
31e40804
105c0554
a0bc0807
08560be7
00000804
40c31016
0824305c
301c6fd2
311c111c
6c0c0000
0c64035c
400614c3
0be4e8bc
4ebc04c3
08560bc0
00000804
201c30c3
211c111c
480c0000
0c44025c
400613c3
0be4e8bc
00000804
50c37016
8c0c616c
0173c006
14c305c3
0bd528bc
0b0d303c
7f327fe5
900cd980
156c96f2
6bd2606c
09e4305c
305c68d2
333c0e04
33c40b0d
d9807f32
0e5606c3
00000804
ff96f016
61c350c3
301c72c3
311c111c
6c0c0000
0c44035c
400615c3
0be522bc
11540007
64ac356c
0d946027
0153840c
14c305c3
0bd528bc
73cc04f2
21946007
97f2900c
111c401c
0000411c
035c700c
15c30c44
e8bc4006
700c0be4
0c44335c
40374006
17c306c3
35c323c3
0be53cbc
1150001c
0000011c
40062806
09d926bc
0f560196
00000804
000620c3
31c32829
31832849
31832809
31832869
31832889
318328a9
00ff331c
00260294
00000804
10fc301c
0000311c
6c0c6c0c
20c30e49
103c0e69
20a7412c
035c1094
10c30119
0121035c
40ac203c
0026323c
fff0133c
fff0323c
00f331a3
fff0213c
0026313c
32a37fe5
f88c033c
00000804
10fc301c
0000311c
6c0c6c0c
05e1035c
00000804
ff961016
326432c3
644c6037
233c6ccb
241c400c
6832ffff
301c23a3
311c88c7
43c30000
0e9424e4
0bb4301c
0000311c
6e2c6c2c
2161235c
341c32c3
69f20020
301c02b3
311c888e
43c30000
0e9424e4
1110301c
0000311c
335c6c0c
4f5c0724
24c30001
01643664
00060053
08560196
00000804
51c33016
10fc301c
0000311c
8c0c6c0c
0bc254bc
00070164
a0272a54
52492894
526912c3
40ac323c
145460a7
0de9345c
10546007
0e546067
3051145c
341c31c3
60070008
245c1154
4ed20b69
07c9345c
301c6bd2
311c111c
6c0c0000
08e4335c
36640026
20260093
0b7d145c
0c560006
00000804
ff96f016
601c40c3
611c0bb4
782c0000
502b0e0c
2249b100
226971c3
43ac313c
0005361c
133c7fe5
2037f90c
138375e9
145c2037
f4890283
62056b80
704f7180
37c3f0cb
6d207e05
6d205489
208770ce
301c1694
311c1110
6c0c0000
0744335c
366414c3
e006746c
000f711c
20063783
0001111c
32e421c3
04332694
3f5c14c3
23c30001
0bc284bc
00070164
301c1c94
311c1110
6c0c0000
0464335c
7f5c04c3
17c30001
746c3664
111c2006
3183000f
211c4006
72c30001
059437e4
14c3180c
08e71abc
0f560196
00000804
0736f016
90c350c3
9184202b
1110301c
0000311c
19c36c0c
335c440c
023c07a4
3664fff4
000780c3
a55c2854
78c30293
0413c006
29c3cdf2
31c32889
07c36205
54cb2980
0bcdb4bc
fd0054cb
363c01f3
263c0010
9500180c
153c07c3
243c3e1d
b4bc063e
700b0bcd
363cfd80
63c30010
6ae46364
08c3e014
0f56e076
00000804
01c330c3
27f262d2
00a4001c
0a7762bc
00f31fe6
0300133c
b4bc40c6
00060bcd
00000804
201c30c3
211c10fc
480c0000
13c3080c
b0bc40c6
080408cb
0736f016
40c3fd96
a3c351c3
01649f5c
836482c3
001c06f2
62bc00a5
0d730a77
111c301c
0000311c
4c4c6c0c
31c3280b
680e6025
1110301c
0000311c
335c6c0c
030607a4
70c33664
00077fe6
000942dc
40c615c3
0bcdb4bc
02f9245c
602647f2
02fd345c
b0bc05c3
673c0bc3
06c30060
4800143c
b4bc40c6
32490bcd
326921c3
412c313c
0e9460a7
143c05c3
40c60300
0bcdd2bc
06c307d2
01d0143c
b4bc40c6
383c0bcd
383c408c
7cce41ac
0063931c
32490b94
326921c3
412c313c
604763d2
62460394
61c60053
1f5c2026
40060006
00252f5c
1ac30006
b2bc29c3
60c30a79
301c0cf2
311c1110
6c0c0000
07c4335c
366407c3
07f37fe6
5489a08c
31c3238b
341c7e05
6e720fff
6026740e
931c744d
1c940063
13c37249
033c7269
03d240ac
14940047
42725469
3f5c40b7
746d0041
433c788c
04c30100
40862006
0bcea4bc
300d3dc6
548d4086
388c4086
033c6880
17c30100
b4bc41c6
06c30bcd
0a8736bc
1110301c
0000311c
335c6c0c
07c307c4
60063664
039603c3
0f56e076
00000804
fc963016
50c340c3
37540007
105c2006
105c02dd
205c02e5
12c30161
0169205c
40ac323c
0171105c
81ac313c
0179205c
c1ac523c
babc0106
00f70bce
00613f5c
0165345c
420b203c
2f5c40b7
245c0041
103c016d
2077440b
00211f5c
0175145c
583220c3
3f5c4037
345c0001
05f2017d
0088001c
0a7762bc
049605c3
08040c56
f096f016
61c370c3
43c352c3
e2dc2007
40070009
000992dc
20072697
000952dc
111c301c
0000311c
4c4c6c0c
31c3286b
686e6025
01400f3c
45862006
0891b0bc
2f5c4026
655700a5
0034233c
3f5c4137
3f5c0081
85d200ad
40bc04c3
04d20bc2
1f5c2046
2f5c00a5
353c00a1
60f7212c
00613f5c
00a53f5c
02e9165c
165c21c3
313c02f1
68d2412c
0f3c87d2
14c30360
b4bc40c6
46970bcd
640732c3
0f3c24b4
26570160
0bcdb4bc
03411f5c
01e51f5c
00a92f5c
500632c3
60b732a3
00413f5c
00ad3f5c
1f5c2026
40060006
00252f5c
1f3c0006
45860140
b2bc30c3
40c30a79
06930bf2
0b84301c
0000311c
001c6c0c
3664220f
a08c0573
744d6606
21c33a49
313c3a69
60a7412c
07c30c94
f7cc101c
0017111c
d2bc4066
03f20bcd
74ed6026
31c3338b
341c7e05
6e720fff
4086740e
01d5245c
365c6026
200602cd
02d5165c
36bc04c3
00060a87
1fe60053
0f561096
00000804
fc96f016
301c60c3
311c111c
6c0c0000
282b4c4c
602531c3
70c3682e
42890cd2
42a912c3
40ac323c
313c22c9
42e981ac
c1ac723c
00805f3c
200605c3
b0bc4106
301c0891
311c111c
6c0c0000
0c04435c
15c30c6c
46644106
416440c3
05c9165c
165c21c3
313c05d1
6287412c
165c3e94
21c309d9
09e1165c
412c313c
09e9265c
81ac323c
09f1165c
c1ac213c
40074077
2f5c2c94
265c0021
32c305cd
05d5365c
7f2ce9d2
0200331c
375c0594
60070ba4
5a491c94
5a6912c3
40ac323c
08946047
0c84375c
211c4006
32830002
301c6ef2
311c111c
6c0c0000
20066ccc
01c32037
36c323c3
0be53cbc
049604c3
08040f56
0c0c616c
634c0173
0200341c
305c66d2
63f20e04
00730026
16f2000c
00000804
301cfe96
311c1398
6c0c0000
07d46047
20e4305c
0fc364d2
0bcd92bc
08040296
60c3f016
305c71c3
a00620e4
13546007
353c01b3
265c0187
8d0020e4
17c304c3
d2bc40c6
08d20bcd
365ca025
23c32104
f01452e4
04c38006
08040f56
205c4006
305c2147
6ad22124
0bc5febc
606c07d2
606f6025
92bc0205
08040bcd
0136f016
41c350c3
101c01c3
111cf204
54bc0050
00070bc0
04c35454
f204101c
0050111c
0bc168bc
000760c3
153c4a54
40260140
0bcf9abc
004770c3
e0060554
02940027
06c370c3
0bcf06bc
0530843c
18c305c3
0bc5febc
0cd260c3
37e4604c
e04f3054
2d54e007
16c305c3
0bd2febc
301c0513
311c1110
6c0c0000
2104255c
0804335c
20e4055c
0010123c
36644306
17540007
20e7055c
2104255c
0187323c
323c8180
355c0010
04c32107
430616c3
0bcea4bc
18c304c3
b4bc40c6
f04f0bcd
0f568076
00000804
60c37016
800651c3
740c0113
133c06c3
2cbc4a1d
80250bc6
32c3542c
f61443e4
eebc06c3
0e560bc5
00000804
0136f016
6007624c
305c2e94
60a707e4
60c32ab4
5a4e563c
0140703c
111c801c
0000811c
05c303d3
f204101c
0050111c
0bc89ebc
000740c3
7ebc1354
20c30bcf
04c30cf2
9abc17c3
07f20bcf
680c28c3
08c4335c
366404c3
06bc04c3
b40c0bcf
e29456e4
0f568076
00000804
1f36f016
a1c350c3
0800023c
0bea00bc
000740c3
0ac35454
f204101c
0050111c
0bc89ebc
80c390c3
301c0ad2
311c111c
6c0c0000
08a4335c
80c33664
573c75c3
ba3c5a4e
c01c0200
c11c111c
06330000
2e545ae4
101c05c3
111cf204
9ebc0050
40c30bc8
24540007
0bcf7ebc
1d540007
680c2cc3
08a4335c
366404c3
0bc360c3
0200153c
d2bc40c6
0fd20bcd
68d238c3
08c3c7d2
420616c3
0bcdd2bc
04c306d2
0bcf06bc
01138026
06bc04c3
b40c0bcf
cf9457e4
09c38006
0bcf06bc
f87604c3
08040f56
0136f016
61c380c3
413c72c3
04c30800
0bea00bc
10540007
101c07c3
111cf204
9ebc0050
50c30bc8
21540007
0bcf7ebc
27940007
04c30393
0be9e4bc
000750c3
07c31654
f204101c
0050111c
0bc89ebc
0dd250c3
0140183c
9abc4026
00070bcf
28c31094
0964325c
0bd46047
6bd2798c
0180063c
0200173c
d2bc40c6
03f20bcd
00538026
05c38006
0bcf06bc
807604c3
08040f56
60c37016
02c351c3
341c674c
60070200
101c3554
111cf204
9ebc0050
40c30bc8
0080521c
00bc05c3
0ad20bea
28548007
7ebc04c3
50c30bcf
1b940007
05c30293
0be9e4bc
14540007
1a548007
163c04c3
40260140
0bcf9abc
0bf250c3
0964365c
07d46047
06bc04c3
05c30bcf
86d20153
06bc04c3
00260bcf
1fe60093
00060053
08040e56
403c1016
04c30800
0bea00bc
04c306f2
0be9e4bc
02d26046
03c36026
08040856
000620c3
31c32829
31a32849
31a32809
31a32869
31a32889
31a328a9
002662f2
00000804
0804002c
0804004c
0bc7eebc
00000804
200c21c3
082f280f
442f200c
0804400f
f4bc002c
08040bc7
602c200c
602c642f
60062c0f
602f600f
00000804
00000804
600c0dd2
600f7fe5
301c69f2
311c1110
6c0c0000
07c4335c
08043664
0644205c
205c4025
40060647
06a7205c
00000804
20c33016
426441c3
0084021c
21806bcc
a0290153
404525c3
08d423e4
34e46009
01000654
60276420
0006f5d4
08040c56
30c37016
021c51c3
4fcc0084
03738100
313c2029
32e40020
600919d4
00dd331c
20670f94
60690d35
c0497012
c1ac363c
32a340a9
363cc089
53e441ac
313c0854
01800020
40275020
0006e4d4
08040e56
51c37016
400743ec
303c2454
23cc0840
81000c80
20290373
0020313c
19d432e4
331c6009
0f9400dd
0d352067
70126069
363cc049
40a9c1ac
c08932a3
41ac363c
085453e4
0020313c
50200180
e4d44027
0e560006
00000804
41c33016
28d252c3
22bc12c3
14c30bcf
b4bc25c3
0c560bcd
00000804
0136f016
81c350c3
40bc03cc
60c30bcf
35540007
0840453c
f00017cc
54c30493
009e253c
0020323c
20d431e4
331c7009
159400dd
13354067
70127069
303c1049
30a9c1ac
108931a3
41ac303c
079483e4
143c06c3
5f850060
0bc890bc
32c35409
91806045
20273e20
06c3dbd4
0bc7ecbc
05f240c3
06bc06c3
64c30bcf
807606c3
08040f56
50c33016
31c341c3
29cf033c
053c14ef
13c30200
b4bc40c6
502c0bcd
708b568f
02a6355c
055c10ab
506c02b6
708c56cf
10ec76ef
70cc170f
572f50ac
053c774f
92bc06c0
710c0bcd
03e8101c
2310141d
0d20776c
710c176f
3310341d
128d133c
21e4578c
303c0a15
776ffff0
4240001c
000f011c
778f6800
6ca0778c
0c56778f
00000804
0136f016
61c370c3
2d542007
2006044c
01930af2
7e8c582c
1a1d423c
35e454c3
20250554
f71410e4
7b2c0413
1b546007
02c0873c
a00646c3
106c0233
13540007
4007508c
7e6c1054
21e413c3
18c30594
0bcdd2bc
a02508d2
5b2c8105
53e432c3
0073ed14
00530026
80760006
08040f56
51c37016
8c0c616c
02c0613c
108c0213
50ac0dd2
366c4bd2
23e431c3
16c30794
0bcdd2bc
002603f2
900c0093
04c391f2
08040e56
50c33016
228c41c3
275441e4
526c2dd2
03c3666c
239420e4
02c0043c
d2bc2585
00070bcd
84051c94
dabc04c3
00070bc7
04c31694
0380153c
d2bc40c6
0dd20bcd
153c04c3
40c603e0
0bcdd2bc
0b0d303c
033c7fe5
0093f88c
00530026
0c560006
00000804
0336f016
81c390c3
101c01c3
111cf204
9ebc0050
60c30bc8
000740c3
7ebc3754
50c30bcf
0bf2e026
193c06c3
27c30140
0bcf9abc
75c340c3
25540007
616c09c3
583c8c0c
03b302c0
341c734c
60070200
50ac1754
18c34bd2
03c3666c
109420e4
15c3108c
0bcdd2bc
043c0bf2
e4d20800
0bea00bc
e4bc0073
40c30be9
900c0093
e3948007
06bc06c3
04c30bcf
0f56c076
00000804
fd96f016
41c330c3
46474077
40573454
264712c3
12c308b4
2d542027
260712c3
05331294
32c34057
f201201c
0050211c
0b5432e4
13c36057
f204301c
0050311c
0c5413e4
0df38006
3cbc2057
70c30bc8
205704c3
0bc054bc
205703d3
0bc89ebc
04c350c3
68bc2057
60c30bc1
a00775c3
03531794
00211f5c
03c320b7
00412f5c
24bc12c3
70c30bc8
3f5c04c3
13c30041
0a812cbc
37c340c3
1b94e007
05c303b3
0bc7f0bc
46c370c3
06c3c5d2
0bc7f0bc
35c340c3
05c3a5d2
0bc7ecbc
06c330c3
1454c007
603706c3
0bc7ecbc
01d36017
31c33c29
85f26045
54c304c3
00d364c3
02c35029
a0060045
e2d265c3
373c8cf2
233c0b0d
343cfff0
7fe50b0d
433c3283
0173f88c
089430e4
14c307c3
d2bc23c3
80260bcd
800602d2
06bc05c3
06c30bcf
0bcf06bc
039604c3
08040f56
50c37016
04ab61c3
055c20c3
200302b3
768c8006
01c3242c
025430e4
770c8026
01c338ec
025430e4
323c8172
62d20104
323c8272
62d20024
57cc8372
31c3392c
099423e4
0840053c
05c0163c
0bcdd2bc
2a540007
05c38872
201c16c3
211cf201
f0bc0050
02f20bc9
05c38472
460616c3
0bc9f0bc
857202f2
16c305c3
f204201c
0050211c
0bc9f0bc
867202f2
16c305c3
f0bc4026
07d20bc9
16c305c3
f0bc4646
02f20bc9
04c38772
08040e56
60c37016
52c341c3
0014313c
288c64d2
0be7a6bc
0024343c
06c365d2
a8bc348c
343c0be7
65d20044
348c06c3
0be7aabc
0084343c
06c365d2
acbc348c
343c0be7
65d20104
348c06c3
0be7aebc
0204343c
06c365d2
b0bc348c
343c0be7
65d20404
348c06c3
0be7b2bc
1004343c
06c365d2
b4bc348c
343c0be7
65d20804
348c06c3
0be7b6bc
08040e56
0736f016
41c370c3
01c352c3
86bc12c3
90c30bca
30af2006
0644275c
04c350cf
e0bc15c3
04c30bc8
0bc800bc
101c04c3
111c9a09
3cbc506f
0ad20bc8
101c05c3
111c9a09
54bc506f
00070bc0
754c5254
4c80352c
33cc73ec
32e46c80
043c0c14
153c0840
b4bc05c0
352c0bcd
554c33cf
07f353ef
043c1070
00bc0080
301c0bc8
311c1110
4c0c0000
354c752c
225c6c80
04c307e4
0840133c
60c32664
24540007
06a4075c
01934006
100c123c
0684375c
640c2580
039434e4
0093c40f
20e44025
7e8cf414
029434e4
754cde8f
0840063c
05c0153c
4e00952c
0bcdb4bc
3bcf352c
5bef554c
08c346c3
0080143c
0bc7f4bc
0b40073c
fcbc14c3
07c30bc7
24c319c3
0bcadcbc
e07604c3
08040f56
0136f016
81c340c3
63c372c3
0bc088bc
19540007
453c54c3
02735a4e
0200043c
40c618c3
0bcdd2bc
726c0bf2
089436e4
02c0043c
26c317c3
0bcdd2bc
900c05d2
ed9445e4
04c38006
0f568076
00000804
0136f016
51c340c3
0684105c
1f542007
06a4605c
03330006
100c703c
0a1d313c
0010203c
109435e4
78204212
07806212
233c2500
bebcffc0
345c0bcd
7fe506a4
06a7345c
02c30093
e71406e4
00bc05c3
053c0bc8
00bc0080
345c0bc8
7fe50624
0627345c
111c301c
0000311c
335c6c0c
04c30884
0200153c
3664548c
0cbc17ac
301c0bc8
311c1110
6c0c0000
07c4335c
366405c3
0f568076
00000804
0136f016
81c350c3
021c42c3
92bc00e0
08c30bcd
600c04d2
30946007
2e548007
463c65c3
f00c5a4e
05c304f3
74bc14c3
00070bc9
04c31f94
22bc18c3
00070bc9
70cc1954
0644155c
32e421c3
70ac0434
70af6025
70ac556c
0924025c
31e410c3
05c30914
201c14c3
211cf7d0
cebc0017
47c30bcb
46e4fc0c
8076d994
08040f56
60c3f016
453c50c3
03135a4e
14c306c3
0bc95abc
11940007
14c306c3
0bc9a6bc
0bf270c3
14c306c3
f804201c
0017211c
0bcbcebc
00b307c3
45e4900c
1fe6e894
08040f56
60c3f016
0bcc5cbc
600730c3
56c31954
5a4e453c
06c30253
74bc14c3
70c30bc9
06c30bf2
201c14c3
211cf7ec
cebc0017
07c30bcb
900c00b3
ee9445e4
0f561fe6
00000804
0136f016
81c360c3
43c372c3
114c6d2c
033c6c00
babc0840
50c30bce
4b540007
0664365c
6025608f
0667365c
0644165c
14c320cf
0bc8e0bc
02c0053c
27c318c3
0bcdb4bc
512cf66f
714c57cf
714c77ef
0840053c
05c0143c
4f80f12c
0bcdb4bc
0624365c
0010233c
035c796c
10c308e4
0b3521e4
7ebc06c3
07d20bcc
265c796c
40250624
08e7235c
0b40063c
fcbc15c3
063c0bc7
153c0bc0
fcbc0080
365c0bc7
60250624
0627365c
153c06c3
548c0200
0be7a4bc
807605c3
08040f56
0136f016
71c350c3
200601c3
0a812cbc
000740c3
60c37a54
009e363c
75b46407
101c07c3
111c9a09
54bc506f
05f20bc0
1884355c
0d336fd2
40e75809
043c0b94
101c0020
111cf7e4
d2bc0017
00070bcd
80455c54
173c05c3
24c30530
a6bc7809
10c30bcb
05c309f2
580914c3
a0bc37c3
60c30bcc
05c302d3
20bc27c3
60c30bcb
0684155c
055c2ed2
400606a4
323c0113
8581100c
68e484c3
40253854
f81420e4
3354c007
0161475c
0405465c
06c4255c
06a4355c
1f1432e4
43d28306
080c423c
1110301c
0000311c
335c6c0c
055c0804
14c30684
36644086
301c0af2
311c0b84
6c0c0000
220e001c
01f33664
0687055c
06c7455c
0684255c
355c48d2
623c06a4
60253b9d
06a7355c
0f568076
00000804
10f0301c
0000311c
201c6c0c
211c86a0
033c0001
0804228d
40c31016
0bcd86bc
4e24102f
301cf524
311c10f4
6c0c0000
323c700f
62d24004
0006f324
08040856
40c31016
0bcd86bc
301c102f
311c10f4
6c0c0000
0006700f
08040856
60061016
85a200b3
602581a1
5cf25fe5
08040856
50c37016
01e442c3
b4bc0434
01530bcd
26004100
00936006
09a105a2
7fe59fe5
05c39cf2
08040e56
50c37016
12c341c3
45f26006
60250153
075413e4
11a255a2
fa5420e4
00530820
0e560006
00000804
005330c3
40090025
01a05ef2
00000804
50c37016
000740c3
e6bc1454
603c0bcd
301c0010
311c1110
6c0c0000
07a4335c
366406c3
05d240c3
26c315c3
0bcdb4bc
0e5604c3
00000804
00d330c3
039401e4
009303c3
0c086025
08041af2
20c31016
005330c3
0c096025
033c1ef2
00b3fff0
31e46008
1fe50554
fb3402e4
08560006
00000804
40c33016
400601c3
402500b3
03c363f2
710200f3
31e42102
03c3f954
01a031c3
08040c56
0bce28bc
00000804
50c37016
12c341c3
48f26006
03f201f3
015330c3
13e46025
15820954
02e45182
30c3f754
0c2002c3
00060053
08040e56
0bce3ebc
00000804
40c31016
12c301c3
00f34006
71216122
40256102
62d23fe5
04c33af2
08040856
fe961016
01c330c3
12544007
01534077
008f203c
4f5c4037
8c0d0001
10544007
40576025
9fe542c3
93f28077
303c00b3
7ef2008f
2f5c00b3
4c0d0021
31e3ff33
02960180
08040856
40c37016
01c351c3
0bcde6bc
015360c3
15c304c3
3ebc26c3
03f20bce
009304c3
10088025
0e5616f2
00000804
ff961016
203740c3
30c312c3
49f24017
08cb9cbc
2f5c00f3
233c0001
3fe500df
04c33bf2
08560196
00000804
50c33016
1110301c
0000311c
335c6c0c
366407a4
05d240c3
25c32006
0bcea4bc
0c5604c3
00000804
30c33016
501c41c3
511c111c
540c0000
13c3080c
f6bc24c3
40c30b1b
1e540007
10fc301c
0000311c
6c0c6c0c
0bc1035c
035c10c3
203c0bc9
135c40ac
213c0bd1
035c812c
303c0bd9
6027c12c
80060354
740c00b3
0864335c
04c33664
08040c56
0804002c
0804004c
0bcf00bc
00000804
40c31016
17540007
341c606c
6ad20001
1110301c
0000311c
335c6c0c
004c07c4
301c3664
311c1110
6c0c0000
07c4335c
366404c3
08040856
40c3f016
02bc51c3
70c30bcf
febc04c3
60c30bce
7480302c
500c702f
31e412c3
301c0b35
311c111c
6c0c0000
0cc4335c
15c304c3
1f003664
08040f56
40c31016
babc0205
05d20bce
433c30c3
604f087f
08040856
ff961016
0484305c
18546007
20072c09
020c1554
00076026
40061254
14c38029
343c8009
316440ac
02946087
423c4026
80370016
00013f5c
60060053
019603c3
08040856
83961016
88bc1fc3
30c30bd2
30e40006
0fc30474
0bcf4cbc
08567d96
00000804
1fc38396
0bd288bc
13740007
60076917
4c091054
64174ed2
00066cd2
21c32c29
313c2c09
3164412c
04946087
00530026
7d960006
00000804
0136f016
40c38196
62c371c3
1f600f3c
f824101c
0017111c
e6bc40c6
04c308cb
88bc1fc3
00070bd2
60572874
c5d266f2
4cbc0fc3
04530bcf
a0069097
0006801c
1f606f3c
14948007
04c30313
40c617c3
0bcdd2bc
004603f2
04c30233
40c616c3
0bcdd2bc
002603f2
80c50133
70d7a025
3380141d
ea1453e4
7f960006
0f568076
00000804
0804002c
0804004c
40c37016
60062364
2e354047
56c3c449
363cc409
a42982ac
41ac353c
372a331c
301c0d94
311c111c
6c0c0000
0844335c
5fa52065
30c33664
231c02f3
13b40400
0f84005c
0fb40127
0680303c
3b9d143c
0720303c
3b9d243c
0010303c
0f87345c
00536006
03c37fe6
08040e56
42c31016
23c31364
131c2364
e2dc1028
131c001b
b5dc1028
131c0008
42dc1014
131c0018
42b41014
1009131c
0014f2dc
1009131c
131c1eb4
92dc1003
131c0019
0ab41003
1001131c
002432dc
1002131c
002464dc
131c26d3
72dc1005
131c0015
c0dc1005
131c0010
94dc1008
22b30023
100f131c
001812dc
100f131c
131c0ab4
62dc100d
131c0010
94dc100e
3a530022
1011131c
001b92dc
1011131c
000f40dc
1012131c
0021c4dc
131c22d3
42dc1020
131c0017
1eb41020
1017131c
0014e2dc
1017131c
131c0ab4
32dc1015
131c0013
54dc1016
27930020
101a131c
000bb2dc
101e131c
0013f2dc
1018131c
001f84dc
131c3393
92dc1023
131c0017
0ab41023
1021131c
0016d2dc
1022131c
001e84dc
131c1393
52dc1026
131c0013
25dc1026
131c001a
b4dc1024
2c93001d
1044131c
000e72dc
1044131c
131c42b4
c2dc103c
131c000b
1eb4103c
1032131c
001642dc
1032131c
131c0ab4
22dc102c
131c000c
d4dc102d
18f3001b
103a131c
0012d2dc
103a131c
0012f5dc
1039131c
001b04dc
131c0dd3
a2dc103f
131c000d
0ab4103f
103d131c
000bf2dc
103e131c
001a04dc
131c17d3
a2dc1041
131c0010
b0dc1041
131c000c
34dc1042
24330019
1053131c
131c7154
1cb41053
1048131c
131c5254
0ab41048
1045131c
0013e2dc
1047131c
0017e4dc
131c0833
2a54104a
104a131c
001690dc
104d131c
001724dc
131c27b3
52dc1059
131c0013
0db41059
1055131c
0014c2dc
1055131c
131c4a14
f4dc1057
25f30015
1062131c
000c32dc
106a131c
0012d2dc
1061131c
001524dc
40271673
0014c4dc
2973800f
74dc4027
804f0014
420728d3
001424dc
2833806f
d4dc4207
808f0013
42072793
001384dc
26f380cf
34dc4207
80af0013
40472653
0012e4dc
25b380ef
94dc4047
810f0012
40272513
001244dc
2473812f
f4dc4047
814f0011
404723d3
0011a4dc
2333816f
54dc4107
818f0011
40272293
001104dc
21f381af
b4dc4047
81cf0010
40472153
001064dc
20b381ef
14dc4047
820f0010
323c2013
3364fda0
95dc6207
405c000f
205c08c7
1eb308e7
14dc4087
822f000f
40271e13
000ec4dc
1d73824f
74dc4107
826f000e
44071cd3
000e24dc
1c33828f
d4dc4407
82af000d
44071b93
000d84dc
1af382cf
34dc4407
82ef000d
42071a53
000ce4dc
19b3830f
94dc4207
832f000c
42071913
000c44dc
1873834f
f4dc4207
836f000b
410717d3
000ba4dc
1733838f
54dc4047
83af000b
40471693
000b04dc
15f383cf
b4dc4027
83ef000a
40271553
000a64dc
0407405c
40c71493
000a04dc
0427405c
402713d3
0009a4dc
0447405c
40271313
000944dc
0467405c
40271253
0008e4dc
0487405c
40271193
000884dc
04a7405c
402710d3
000824dc
04c7405c
405c1013
205c0587
0f7305a7
05c7405c
05e7205c
405c0ed3
205c0607
0e330627
0647405c
0667205c
44070d93
405c6ab4
205c0687
0cb306a7
f420323c
60473364
405c60b4
205c06c7
0b7306e7
0707405c
0727205c
105c0ad3
21270b84
313c52b4
403c0480
313c3b9d
203c0520
313c3b9d
305c0010
08b30b87
43b44407
0747405c
0767205c
405c07d3
205c0787
073307a7
07c7405c
07e7205c
405c0693
205c0807
05f30827
2b944027
04e7405c
41070553
105c2694
21270ce4
313c24b4
403c05d0
313c3b9d
305c0010
03730ce7
0080231c
323c16b4
60070074
405c1294
205c0887
03c308a7
14c301f3
0bcfe0bc
09150007
404700d3
405c0494
00730567
00531fe6
08560006
00000804
0336f016
91c340c3
200601c3
01f4201c
0bcea4bc
debc04c3
50c30bcf
dcbc04c3
85c30bcf
00068084
28c30733
60676aa0
25c338f4
009e323c
613c3409
35c341ac
011e433c
2c298812
733c41a3
38c30020
41e42fa0
641c0af4
631cff00
21541000
1027031c
03331e94
36a334c3
05c36cf2
00b323c3
00256089
402564f2
fb7421e4
115421e4
16c309c3
34c327c3
0bd016bc
07740007
06c35e00
58e452c3
0073c714
00531fe6
c0760006
08040f56
60c3f016
0904005c
265c4006
52c30907
1110701c
0000711c
606c0173
021553e4
800c53c3
335c7c0c
366407c4
16f204c3
0924365c
365c6e80
0f560927
00000804
60c3f016
000771c3
20072454
405c2254
a0060904
043c0393
17c30040
d2bc40c6
00070bcd
700c1294
365ca4f2
00530907
301c740f
311c1110
6c0c0000
07c4335c
366404c3
00d30006
900c54c3
e4948007
0f561fe6
00000804
51c33016
23f202d2
01b38006
0904405c
043c0133
15c30040
d2bc40c6
03d20bcd
98f2900c
0c5604c3
00000804
50c37016
26540007
601c8006
611c1110
01330000
4a1d003c
780c05d2
07c4335c
80253664
542c140c
43e432c3
09d2f414
1110301c
0000311c
335c6c0c
366407c4
1110301c
0000311c
335c6c0c
05c307c4
0e563664
00000804
000620c3
31c32829
31a32849
31a32809
31a32869
31a32889
31a328a9
002662f2
00000804
0804002c
0804004c
40a1041c
002602d2
00000804
0542041c
002602d2
00000804
40c31016
0bd382bc
07f26026
88bc04c3
02d20bd3
30c30026
085603c3
00000804
40c31016
0bd38ebc
03f26026
090b343c
085603c3
00000804
111c301c
0000311c
335c6c0c
03ac0824
08043664
305c20c3
6c6c0744
63d21fe6
36640bac
00000804
fa96f016
61c350c3
13c372c3
0744205c
1fe6688c
17546007
355c6006
77ac08e7
22d72037
23172077
235720b7
239720f7
23d72137
888c2177
01a0053c
26c313c3
466437c3
0f560696
00000804
305c20c3
6dec0744
63d21fe6
36640bac
00000804
0744305c
63d26e0c
366403ac
00000804
305c20c3
6e8c0744
63d203c3
36640bac
00000804
50c33016
0744005c
04c382ac
17ac83d2
0c564664
00000804
00000804
00000804
08040006
00000804
0136f016
80c3fb96
61c371c3
1540513c
04c38006
0ca4265c
16544007
175c34c3
31030d24
0b0d333c
7f327fe5
60066037
60b76077
4137a0f7
202608c3
34c323c3
0bd3bebc
80250026
a205c085
e3948087
80760596
08040f56
60c3f016
22a4305c
29546007
701ca006
711c1110
02530000
0387453c
42007c0c
07c4335c
3664084c
365c5c0c
6e0022a4
07c4225c
26640c8c
365ca025
065c22c3
53e422a4
301cea74
311c1110
6c0c0000
07c4335c
60063664
22a7365c
08040f56
fb967016
61c350c3
08e4405c
58948007
80778037
80f780b7
14c38137
34c324c3
0bd3bebc
80778037
80f780b7
05c38137
24c314c3
bebc6026
80370bd3
80b78077
813780f7
14c305c3
604624c3
0bd3bebc
80778037
80f780b7
05c38137
24c314c3
bebc6066
80370bd3
80b78077
813780f7
14c305c3
608624c3
0bd3bebc
80778037
80f780b7
05c38137
24c314c3
bebc60a6
c0070bd3
80371254
80b78077
813780f7
14c305c3
34c326c3
0bd3bebc
16c305c3
602624c3
0bd400bc
355c6026
059608e7
08040e56
00000804
00000804
008730c3
00871154
000608d4
0c546027
60470026
01130894
62070066
00a60554
02546807
08040046
040760a6
04072b54
604611d4
26540087
05d40087
00276006
04132094
01076066
60861d54
19940207
61060333
0100031c
031c1554
09d40100
080760c6
60e60f54
0080031c
01530a94
031c6126
06540200
031c30c3
02544000
03c36026
00000804
08040006
616c20c3
00266cac
05546047
0a04325c
0c8b033c
00000804
41c3f016
30542007
0e04315c
2c946007
305c07d2
64d22284
0a24005c
1fe60053
400614c3
0104603c
0024503c
0001041c
0ca4315c
60a76cd2
09f20394
61a702b3
a5f20394
62070233
ced20f94
20854025
ef944087
88bc134c
08d20bd3
66f272ac
72ec03c3
002664f2
00060053
08040f56
600629d2
10a7315c
10c7315c
315c43d2
08041087
50c3f016
62c371c3
0464305c
1b546007
20078006
02f31394
0247343c
0464255c
650c2d00
62e423c3
07c30894
d2bc26c3
03f20bcd
01130026
355c8025
23c30484
eb1442e4
0f560006
00000804
50c37016
305c61c3
80060424
02736ff2
0067343c
0424255c
16c30d00
d2bc40c6
03f20bcd
01130026
355c8025
23c30444
ef1442e4
0e560006
00000804
fe963016
a007a26c
774c3354
0200331c
355c2f54
233c1084
255c0010
355c1087
69d20fc4
19c4305c
22946007
1a04305c
1e946007
012c401c
0eb44647
42878f06
87860bb4
08b44147
40a783c6
828605b4
02b44027
0fc38146
0bcd92bc
70802017
10a4255c
31e412c3
355c03f4
029610a7
08040c56
9ebc03ac
08040bc3
0336f016
50c3f696
00201f3c
0bd3b4bc
000760c3
05c36274
02201f3c
0bd5e8bc
5b740007
60ac156c
0000801c
355c65f2
833c0a04
800c090b
02207f3c
00209f3c
05c30933
28bc14c3
00070bd5
70ac1894
62e423c3
09c30794
26c3308c
0bcdd2bc
38c303d2
718c6cd2
38546007
143c07c3
40c60180
0bcdd2bc
30540007
14c305c3
0bd528bc
15940007
341c734c
60070200
708c1054
70ac63d2
718c6cf2
1e546007
143c07c3
40c60180
0bcdd2bc
16540007
14c305c3
0bd528bc
718c0cf2
70ac6ad2
07c368f2
0180143c
d2bc40c6
06d20bcd
8007900c
0053b794
04c38006
c0760a96
08040f56
0736f016
60c3ee96
52c391c3
2007a3c3
001852dc
101c01c3
111cf201
3cbc0050
40c30bc8
260609c3
0bc824bc
000770c3
778c1e54
0002341c
19546007
12c34029
2f3c2045
c2bc0280
00070be0
772c1094
31832317
770c6cd2
328342d7
774c68d2
31832357
0002801c
41946007
22dc8007
778c0015
0001341c
c2dc6007
04c30014
12c35029
2f3c2045
c2bc0280
00070be0
001414dc
2317772c
60073183
0013b2dc
42d7770c
60073283
001352dc
2357774c
801c3183
60070001
25931a94
19c304c3
a4bc4406
972c0bce
374c170c
0e84355c
62f24406
833729c3
237702f7
80064477
00b374c3
01448f5c
79c349c3
065c1b51
20660784
6abc28c3
778c0beb
0784065c
233c2106
6abc084b
29c30beb
7aac44f2
1b946007
0784065c
84d224c3
23c37029
14c34045
0bebe6bc
44dc0007
065c000f
27c30784
3c29e4d2
404521c3
babc17c3
00070beb
000e74dc
6317572c
323c2383
22060104
10946007
0404323c
480663d2
323c0273
64d20084
7b0f6106
323c01d3
64d20044
3b0f2086
323c0113
60070024
000c92dc
5b0f4046
62d7570c
323c2383
22060104
13946007
0404323c
480664d2
01d35aef
0084323c
610664d2
01137aef
0014323c
e2dc6007
2026000a
574c3aef
23836357
0204323c
60072406
323c1194
63d20404
04b34806
0804323c
301c64d2
02730080
1004323c
101c65d2
3b2f0100
32c30333
4000341c
201c64d2
02334000
0014323c
602664d2
01937b2f
0024323c
60072046
323ced94
60070104
42067b54
065c5b2f
20c60784
6abc5b2c
065c0beb
20860784
6abc5aec
065c0beb
20a60784
6abc5b0c
44570beb
0e84355c
04946067
335c796c
65d20ea4
01c13f5c
62f26732
323c4006
64d20204
5b6f4406
7b6f0053
0784065c
5b6c20e6
0beb6abc
0784065c
0e84255c
04944067
235c796c
21260ea4
0beb6abc
0784065c
46971ac3
0beec2bc
38940007
88bc174c
40c30bd3
0784065c
2c548007
0340153c
4ebc4406
19c30bec
2a542007
6007758c
f4ac2754
2494e007
000716cc
301c2154
311c111c
6c0c0000
5f3c466c
a0370080
20772406
0804435c
02c0193c
1000301c
065c4664
15c30784
4ebc4406
07c30bec
e6bc03d3
04c30bee
1fe60353
00060313
6b8c02d3
084b333c
0010833c
111c301c
0000311c
4f3c6c0c
335c0280
12c307e4
366424c3
38dc0007
d7b3ffed
e0761296
08040f56
40c37016
605c51c3
206707e4
20062754
0bc1aabc
2294a127
0844345c
1e546007
326c04c3
60bc4026
40060bd5
0927245c
0847245c
202604c3
0bd3f6bc
345c6006
345c2147
301c2167
311c111c
6c0c0000
07c4335c
366404c3
a5d201b3
0354a0a7
0894a0c7
245c4026
04c30847
f6bc2006
545c0bd3
56e407e7
301c1554
311c111c
6c0c0000
07a4335c
15c304c3
366426c3
07e4345c
03546127
0494c127
9ebc04c3
0e560be7
00000804
0136f016
40c3fa96
005cc26c
200607a4
0bfaa2bc
07a4045c
9abc2006
732c0bfa
03546087
05946207
07a4045c
00932046
07a4045c
94bc2006
0f3c0bfa
20060040
a4bc4286
b32c0bce
1794a107
20772026
40b74006
323c5bec
62d20014
323c20b7
64d20024
61726097
345c60b7
341c0a04
63d20010
60b76006
0d30716c
0dc4765c
82bc05c3
00070bd3
a1071194
353c0f54
333c2006
033c0b0d
303cfff0
133cf88c
20370016
00013f5c
60060053
345c6177
e13707a4
00678f5c
163c03c3
2f3c0800
36bc0040
06960bf8
0f568076
00000804
40c31016
111c301c
0000311c
0cac6c0c
400614c3
0be4e8bc
143c04c3
febc0380
08560bd2
00000804
ff96f016
61c350c3
616c72c3
67f26cac
0a04305c
0010341c
15946007
111c401c
0000411c
0cac700c
400615c3
0be4e8bc
6cac700c
40374006
17c306c3
35c323c3
0be53cbc
0f560196
00000804
0736f016
81c350c3
a3c392c3
07e4305c
153560a7
0c84305c
211c4006
32830001
2b546007
1244305c
27946007
153c01c3
40c60380
0bcdd2bc
1f540007
0c04055c
0bcf06bc
111c301c
0000311c
335c6c0c
09c30784
36641ac3
0c07055c
42dc0007
053c000c
92bc1840
053c0bcd
18c318c0
b4bc40c6
17130bcd
153c08c3
40c60380
0bcdd2bc
0b0d303c
fff0233c
355c5f32
323c0c84
355c0c1b
355c0c87
6ed21244
111c301c
0000311c
435c6c0c
05c30764
29c318c3
46643ac3
972c12f3
42dc8087
355c0009
60070864
355c5494
341c0a04
69d20008
88bc04c3
05d20bd3
07e4355c
47546127
c5d2d66c
0de4365c
41546027
82bc04c3
07f20bd3
05548107
431ce146
02940200
301ce8c6
311c10fc
6c0c0000
235c6c0c
32c32d71
0002341c
eb4662d2
2254c007
6007768c
7b4c1f54
0200341c
1a546007
0800063c
0be9e4bc
14540007
101c168c
111cf204
9ebc0050
40c30bc8
153c08d2
40260140
0bcf9abc
e14602f2
06bc04c3
05c30bcf
400617c3
0bd8d4bc
0864355c
355c6025
758c0867
34946007
1140053c
40c618c3
0bcdb4bc
88bc172c
00070bd3
301c1094
311c111c
6c0c0000
0744435c
07a4055c
29c318c3
46643ac3
1ad40007
eebc05c3
355c0bd3
341c0a04
69f20008
0784055c
29c318c3
90bc3ac3
01530bf5
82bc172c
06d20bd3
07a4055c
b2bc2026
e0760bfa
08040f56
3f36f016
70c3b296
92c3a1c3
2384305c
305c7992
005c2387
06bc0c04
00060bcf
0c07075c
125c29c3
313c0de4
275cffe0
60470a04
323c1db4
60070404
003ec2dc
111c401c
0000411c
335c700c
07c30724
366419c3
0a150007
200607c3
0bd804bc
335c700c
36640704
5e917ad3
323c7a93
64d20204
f2dc2007
301c003c
311c1110
6c0c0000
07a4335c
00b0001c
60c33664
301c09f2
311c0b84
6c0c0000
22aa001c
275c68f3
41f70784
201c2006
a4bc00b0
60060bce
0ac37e2f
47540007
1cbc07c3
80c30bd5
41940007
0380473c
6cbc04c3
50c30bd3
18c304c3
a4bc40c6
073c0bce
1a3c03e0
40c60200
0bcdb4bc
07c3a4f2
0be79cbc
26c60ac3
0bc824bc
06d240c3
503c6029
60270020
a00602b4
111c301c
0000311c
335c6c0c
075c0da4
24c30784
302984d2
404521c3
366414c3
3254a007
111c301c
0000311c
335c6c0c
075c0de4
14c30784
04d33664
688c29c3
68ac64d2
1a946007
4cac7d6c
16944047
634c09c3
0200341c
10546007
0947275c
3e2f2026
111c301c
0000311c
6d6c6c0c
200607c3
366421c3
073c59b3
200603e0
a4bc40c6
401c0bce
411c111c
700c0000
06e4335c
366407c3
6e6c700c
366407c3
6dac700c
0784075c
21c32006
29c33664
341c6b4c
6ed20008
0d84325c
325c6bd2
333c0da4
7fe50b0d
f88c233c
6d2060a6
60260053
83b009c3
22f21cc3
2ac3c3c3
46544007
101c0ac3
111cf201
3cbc0050
07f20bc8
26060ac3
0bc824bc
38540007
8f4c39c3
8ebc04c3
00070bd3
431c3154
25544000
315c19c3
60070d44
7d6c0415
0e84335c
65d24006
638c09c3
084b233c
0784375c
03c34037
2a3c2006
39c30200
0be480bc
301c0cf2
311c111c
6c0c0000
06c4335c
07a4075c
36642026
00c8101c
3f3c3377
60371340
1ac307c3
29c304f3
343c8b4c
60070084
3ac31454
11546007
82bc04c3
0dd20bd3
111c301c
0000311c
6d0c6c0c
19c307c3
00063664
0af31377
9ebc04c3
00070bd3
101c1154
337700c8
13403f3c
07c36037
29c32006
02003f3c
0bd65ebc
4c540007
441c44b3
301c0200
311c111c
80070000
6c0c3c54
0684435c
06a4335c
366409c3
50c34664
13540007
0bd37ebc
031c40c3
0db400c8
05c31377
0bd380bc
0f3c30c3
13c30200
b4bc24c3
00730bcd
73776006
06bc05c3
301c0bcf
311c111c
6c0c0000
07c36d0c
366419c3
07d20ac3
02b3105c
341c31c3
64d20010
5bcf4046
60260073
00067bcf
01131f4f
6d0c6c0c
19c307c3
93773664
7c0c9f4f
60076eac
93571b54
111c301c
0000311c
19c36c0c
0fc4115c
535c2037
07c30664
3f3c1ac3
4e000200
00c8301c
56646e20
04740007
6c007357
60067377
1ba7375c
00070ac3
101c1954
111c9a09
9ebc506f
40c30bc8
d2dc0007
301c0021
311c111c
6c0c0000
0644335c
075c3664
04c31ba7
0bcf06bc
07c341d3
11401f3c
0bd51abc
000750c3
8f5c24f4
4f3c09a4
28c30200
3f5c4dd2
2f3c0101
42c30200
06946607
01091f5c
604531c3
3f3c8980
4e200200
14c31280
bebc2884
73570bcd
73776e80
1f3c04c3
25c31140
0bcdb4bc
23d21ac3
02001a3c
70bc07c3
1eec0bd4
0bd4d6bc
1f0c80c3
0bd4d6bc
5f2cb0c3
0046323c
0b0d333c
433c7fe5
85f2f88c
d4c3a026
0b944107
19c307c3
0bd414bc
d5c3a026
543c04f2
d0c30016
331c7f2c
03940200
0393a006
0e946107
6bec29c3
0003341c
74dc6007
3dc3001b
34dc6007
5dc3001b
620701b3
301c0b94
311c111c
6c0c0000
05c4335c
19c307c3
175c3664
21b707e4
20a607c3
0bd804bc
40072ac3
3a3c1454
782f02c0
784f6a6c
1cbc07c3
04d20bd5
618c09c3
3a3c6ed2
780f0200
268c1ac3
00f3386f
488c29c3
39c3582f
784f6cac
205c09c3
40270de4
618c0c94
7d6c6ad2
60476cac
393c0694
780f0180
0427265c
315c19c3
60270de4
215c0894
40070ea4
786c04f4
586f62f2
02003f3c
135778af
191118cf
1f2c7931
0bd4eabc
3f4c194f
997138ef
225c29c3
598f0de4
6f6c39c3
0ac3788f
0401005c
0565065c
21d74006
0c85215c
16c309c3
1540293c
1940493c
0ca4305c
45af62d2
0ca4305c
0085662f
42052085
f59424e4
005c09c3
1aaf0d24
0a04375c
0008341c
794c6fd2
03546027
0a9460c7
6ecc39c3
09c37b4f
64d262ac
0340393c
bb8f7b6f
315c19c3
60670e84
7d6c0494
0ea4335c
60077acf
0ac31454
24bc2606
0fd20bc8
12c34029
2f3c2045
c2bc1140
07f20be0
341c7257
63d200c0
7acf6046
005c09c3
1bef0fc4
325c5c2c
66d211c4
11e4125c
0407165c
5fe60093
0407265c
331c794c
47944000
21c32197
43944127
0784475c
0c24345c
345c6025
ba3c0c27
843c0200
c01c1880
c11c111c
0cc30000
145c400c
045c15a4
017715c4
0007bf5c
3a3c6077
60b70640
00678f5c
3f5c6106
525c0085
04c30624
00a13f5c
343c23c3
56642700
600c0cc3
0604335c
1bc304c3
1ac33664
472c674c
04c7265c
04e7365c
0c24345c
0507365c
0a40063c
410618c3
08cbb0bc
005c0ac3
065c0401
40060565
215c21d7
07c30c85
aabc16c3
30c30bd3
35e4a006
375c2715
341c0a04
63f24000
0413a026
03e0473c
111c301c
0000311c
335c6c0c
07c305e4
366414c3
15c307c3
0bd804bc
15c304c3
a4bc40c6
301c0bce
311c1110
6c0c0000
07c4335c
366406c3
301c0e53
311c1110
6c0c0000
07c4335c
366406c3
62077f2c
301c1394
311c111c
6c0c0000
05c4335c
19c307c3
07c33664
0bd8c0bc
212607c3
0bd804bc
a8d20333
325c29c3
20a60de4
0e946027
7d6c0193
27866cac
08946027
305c09c3
22860de4
02546027
07c32146
d4bc4006
3dc30bd8
07c36fd2
0e801f3c
0bd3e4bc
6f5709f2
0002341c
07c365d2
14bc19c3
7e6c0bd4
39e46cd2
301c0a54
311c111c
6c0c0000
075c6d2c
366407a4
3e719e6c
07c35e91
6cbc19c3
07c30be6
0bd858bc
21c33e6c
115442e4
9abc07c3
01b30be7
2fe60ac3
0bc824bc
e4dc0007
c333ffde
0004801c
cb53b8c3
fc764e96
08040f56
61c3f016
453c50c3
6026009e
73548007
1e3580a7
70126069
373ce049
20a9c1ac
e08931a3
41ac373c
f201101c
0050111c
37e471c3
60c90d94
0a946027
28f220e9
9409080f
604534c3
31c3682f
78200a93
18f460a7
16358267
70126069
343c8049
e0a9c1ac
208937a3
41ac313c
ac04401c
000f411c
37e474c3
303c0794
688f0060
80c70733
60693735
80497012
c1ac343c
37a3e0a9
313c2089
401c41ac
411cac01
74c3000f
099437e4
0060303c
140968af
7f8530c3
03d368cf
ac03101c
000f111c
34e441c3
303c0994
68ef0060
37c3f409
690f7f85
101c01f3
111cac09
41c3000f
089434e4
0060303c
f409692f
7f8537c3
6006694f
0f5603c3
00000804
0736f016
51c340c3
02c362c3
4c862006
0bcea4bc
858484c3
353ce006
94c3fff0
0d939384
231c5009
069400dd
6a5449e4
60077029
54c36754
009e153c
0020313c
03f430e4
0bd3ffe6
07944607
5409984f
604532c3
09d3786f
079446c7
5409996f
604532c3
08d3798f
079446e7
540999af
604532c3
07d379cf
0c944707
24352087
60277049
99ef0394
604706b3
9a0f3394
4ca70633
22270994
9a2f2d35
32c35409
7a4f6045
4fe704f3
9a6f0794
32c35409
7a8f6045
402703f3
9aaf0794
32c35409
7acf6045
464702f3
9aef0794
32c35409
7b0f6045
231c01f3
0c9400dd
18c304c3
febc26c3
70c30bdd
0c740007
e00603d2
54090133
604532c3
38c39180
00270e20
07c392d4
0f56e076
00000804
f7967016
62c350c3
19dc22e7
3ba60009
4006340d
0a06544d
3e46146d
4026348d
000654ad
54cd14ed
13c30026
0be212bc
000701f7
353c7c54
18320080
1f5c01b7
350d00c1
503241d7
0f5c4177
0c2d00a1
283221d7
2f5c2137
4c4d0081
00e10f5c
20260c6d
45c3358d
243c4006
002606de
12bc16c3
02370be2
59540007
04bc06c3
03f20be2
5394c027
021734c3
00f71832
00611f5c
00de133c
50324217
0f5c40b7
0c2d0041
28322217
2f5c2077
4c4d0021
01010f5c
20260c6d
400630ad
343c50cd
03570070
202710c3
4c0d0394
435700f3
004702c3
20060b94
4a062c0d
1e464c2d
1f5c0c4d
2c6d01a1
43570313
020702c3
20060894
4a062c0d
1e464c2d
fe930c4d
21c32357
4000231c
00061294
28060c0d
52c62c2d
0c6d4c4d
4ea06085
ffe0123c
2f5c2037
542d0001
00530ea0
09961fe6
08040e56
f596f016
62c350c3
e49743c3
1004375c
62f24506
12e442c6
000f10dc
340d2606
546d4006
744d6026
14c30046
0be212bc
00070277
000e32dc
0040353c
383210c3
2f5c21f7
548d00e1
303210c3
2f5c21b7
4c2d00c1
28322257
2f5c2177
4c4d00a1
01211f5c
40262c6d
45c34c8d
343c6006
004604de
12bc16c3
02b70be2
e2dc0007
06c3000b
0be204bc
c02704f2
000b74dc
429734c3
41375832
00811f5c
00de133c
50324297
1f5c40f7
2c2d0061
48324297
1f5c40b7
2c4d0041
01412f5c
60264c6d
200670ad
043c30cd
44170070
602732c3
200d0394
241700f3
404721c3
60060b94
21e6600d
5586202d
3f5c404d
606d0201
241707f3
231c21c3
08944000
600d6006
202d2806
404d52c6
6417fe73
240713c3
40060994
61e6400d
3586602d
4066204d
641704d3
280713c3
40060994
61e6400d
3586602d
4086204d
64170353
131c13c3
09940080
400d4006
602d61e6
204d3586
01b340a6
13c36417
0100131c
40064f94
61e6400d
3586602d
40c6204d
403c406d
375c0040
62371584
201c69d2
42370080
04946047
00c0301c
20066237
04c3302d
01012f5c
015f203c
1004375c
60266fd2
306d600d
1004375c
0040043c
0040133c
b4bc4206
043c0bcd
64570140
15946407
1004775c
e8f2e077
00212f5c
3f5c402d
303c0021
2006015f
41e6200d
7586402d
20c6604d
0085206d
133c62a0
2037ffe0
00012f5c
03c3542d
1fe60053
0f560b96
00000804
fd96f016
305c42c3
505c14c4
605c14e4
205c1504
60471524
40370d94
1544305c
00b76077
14c301c3
36c325c3
0bdf9cbc
40370113
14c301c3
36c325c3
0bdf02bc
0f560396
00000804
40c3f016
62c351c3
600927d2
04946607
0be312bc
04c300d3
26c315c3
0be262bc
08040f56
006930c3
0c0910c3
c0ac203c
213c2c29
0c49812c
412c303c
101c0026
111cac00
21c3000f
345432e4
101c0046
111cac01
21c3000f
2c5432e4
101c0106
111cac02
21c3000f
245432e4
101c0206
111cac04
21c3000f
1c5432e4
101c0086
111cac05
21c3000f
145432e4
101c0406
111cac06
21c3000f
0c5432e4
ac08001c
000f011c
333c3003
7fe50b0d
033c7f32
0804300c
006930c3
0c0910c3
c0ac203c
213c2c29
0c49812c
412c303c
4000001c
9600101c
0040111c
32e421c3
00263554
ac01101c
000f111c
32e421c3
00462d54
ac02101c
000f111c
32e421c3
04062554
ac03101c
000f111c
32e421c3
08061d54
ac04101c
000f111c
32e421c3
001c1554
101c0080
111cac05
21c3000f
0c5432e4
ac06001c
000f011c
333c3003
7fe50b0d
033c7f32
0804400c
006930c3
0c0910c3
c0ac203c
213c2c29
0c49812c
412c303c
101c0026
111cf200
21c30050
245432e4
101c0046
111cf201
21c30050
1c5432e4
101c0106
111cf202
21c30050
145432e4
101c0206
111cf204
21c30050
0c5432e4
f205001c
0050011c
333c3003
7fe50b0d
033c7f32
0804100c
006930c3
0c0910c3
c0ac203c
213c2c29
0c49812c
412c303c
101c0026
111cf201
21c30050
1c5432e4
101c0046
111cf202
21c30050
145432e4
101c0206
111cf200
21c30050
0c5432e4
9600001c
0040011c
333c3003
7fe50b0d
033c7f32
0804700c
01076406
01071154
60a608d4
0c540047
008761a6
01130894
03540207
03940807
00536206
03c36006
00000804
06540207
04540807
01076006
60c60294
080403c3
01076046
01071254
004706d4
00870b54
01130b94
02076066
60c60854
04940807
60260093
60060053
080403c3
03540207
03940807
01130026
0086303c
0b0d333c
033c7fe5
0804f88c
313c20c3
6cd20104
ac04001c
000f011c
46544047
f204001c
0050011c
313c0833
001c0404
011cac08
6007000f
313c3994
6cd20084
ac02001c
000f011c
30544047
f202001c
0050011c
313c0573
6cd20044
ac05001c
000f011c
22544047
f205001c
0050011c
313c03b3
6cd20024
ac01001c
000f011c
14544047
f201001c
0050011c
313c01f3
03c30014
001c6bd2
011cac00
4047000f
001c0554
011cf200
08040050
0136f016
61c350c3
02c342c3
44062006
0bcea4bc
300f2026
502f4106
306f504f
708f6006
70af70cf
c00770ef
0008e2dc
b9dcc0e7
74090008
00dd331c
000884dc
363c5429
23e4ffe0
000824dc
70127469
323c5449
34a9c1ac
548931a3
41ac323c
f201101c
0050111c
32e421c3
34c97094
34e921c3
412c313c
60273164
363c6894
6067ff80
053c0bf4
66bc0080
104f0be1
ff40363c
06d46027
1fa604d3
5ed46007
053c0453
400600c0
6009502f
602913c3
40ac833c
200718c3
763c4c54
383cff20
73e4100c
603c4674
a0060020
66bc06c3
702c0be1
702f30a3
ff85c085
58e4a025
00b3f674
60271f66
07133894
1ff4e027
706f6006
21c33809
813c3829
28c3412c
29544007
383cffc5
73e4100c
563c2474
c0060020
9ebc05c3
706c0be1
706f30a3
ff85a085
68e4c025
00b3f674
e0271f26
02931494
11f4e027
12c35409
323c5429
336440ac
0133708f
01131fe6
00d31fc6
00931f86
00531f46
80760006
08040f56
0336f016
41c360c3
02c352c3
44062006
0bcea4bc
340f2046
542f4206
6026544f
2006746f
34cf348f
440634af
800754ef
000a92dc
69dc8067
7809000a
44dc6607
5829000a
ffe0343c
e4dc23e4
58490009
586912c3
40ac323c
60273164
000954dc
80679f85
c0850df4
d4bc06c3
144f0be0
82dc0407
9f850008
07d48027
1fa60573
96dc8007
04d30008
0040063c
342f2006
32c34009
923c4029
39c341ac
76546007
ffe0843c
100c393c
707483e4
0020703c
942c61c3
d4bc07c3
04a30be0
e085142f
fffc821c
69e4c025
041cf574
06d20020
1f660b33
5e948027
831c0bd3
20f40001
9c09146f
9c2914c3
40ac943c
200719c3
821c4f54
393cfffe
83e4100c
673c4974
40c30020
1cbc06c3
746c0be1
746f30a3
821cc085
8025fffc
f57449e4
1f2600d3
0001831c
06f33794
0001831c
580933f4
582942c3
422c323c
748f3364
ffe0183c
28f42027
0020063c
24c38009
343c8029
74af412c
233c3fc5
12e4200c
80060515
1ee694af
00450313
652014cf
12f46067
d4bc0100
30c30be0
1ec614ef
0b946407
1fe60133
1fc60113
1f8600d3
1f460093
00060053
0f56c076
00000804
3f36f016
a0c3ea96
c2c3b1c3
c85743c3
04449f5c
04648f5c
0484df5c
16c303c3
d2bc40c6
5f3c0bcd
7f3c00c0
00070120
05c30915
40c614c3
0bcdb4bc
16c307c3
05c30113
40c616c3
0bcdb4bc
14c307c3
b4bc40c6
09c30bcd
440618c3
0bcdd2bc
0f3c30c3
4f3c0180
60070380
19c30815
b4bc4406
04c30bcd
00f318c3
440618c3
0bcdb4bc
19c304c3
b4bc4406
5f3c0bcd
301c00c0
311c111c
49970000
10544007
49866c0c
df5c4037
49570027
435c40b7
0ac30e04
2cc31bc3
466435c3
6c0c01f3
40374986
0027df5c
40b74957
05a4435c
1bc30ac3
35c32cc3
16964664
0f56fc76
00000804
03d230c3
1004305c
080403c3
600604d2
1007305c
00000804
71c3f016
53c362c3
02f3800c
043ce8d2
17c30400
d2bc40c6
0ef20bcd
043cc8d2
16c30040
d2bc4206
06f20bcd
526ca8d2
53e432c3
900c0454
e9948007
0f5604c3
00000804
0136f016
51c340c3
83c372c3
0fe4605c
205c4006
28d21007
12c306c3
5ebc25c3
045c0be4
373c1007
33c40b0d
f88c533c
1004245c
a8d249f2
17c306c3
5ebc38c3
045c0be4
345c1007
60071004
61971194
aed26fd2
111c301c
0000311c
335c6c0c
06c30544
27c318c3
045c3664
345c1007
333c1004
7fe50b0d
f90c033c
0f568076
00000804
301c3016
311c1110
6c0c0000
70cc8c6c
1b546007
50cf4006
62d270ec
a00650ef
153c0213
70ac200c
686c4c80
600669d2
70ac686f
4c4c6c80
2c2c0c0c
a0252664
32c3508c
ee7453e4
08040c56
1f36f016
91c3b0c3
201c82c3
211c1110
680c0000
6e24ec6c
f524a3c3
80061c6c
c2c364c3
a0ac03d3
3be4608c
604c1894
045439e4
ffff931c
606c1294
045438e4
ffff831c
83f20c94
0053bc6f
2cc3b0af
335c680c
366407c4
0053c025
05c340c3
e2940007
40043a3c
f32462d2
f87606c3
08040f56
40c33016
1110301c
0000311c
6c6c6c0c
01b30c6c
34e4608c
604c0994
069431e4
32e4606c
00260394
00ac0073
0c5614f2
00000804
0336f016
71c350c3
83c392c3
1110301c
0000311c
cc6c6c0c
07a4335c
36640306
7fe640c3
4c540007
0bcd92bc
6e80700c
702c700f
01336f80
6025700c
101c700f
111cbdc0
6880fff0
502c702f
423f301c
000f311c
21e413c3
1051f0d4
706f61d7
20063091
186c30af
6e240bf2
986ff524
0400341c
23546007
30c3f324
ee240433
b00cf524
200620c3
53e4680c
53e40d74
30300694
83c3682c
067498e4
12c368ac
23c363d2
24f2fe53
986f10af
64ac0093
84af70af
4004373c
f32462d2
03c36006
0f56c076
00000804
fe967016
1110301c
0000311c
ac6c6c0c
6007750c
746c3794
742c64f2
32f46007
0be4c2bc
6007746c
0fc32b54
0bcd92bc
f5240e24
946c2017
4026700c
0b7413e4
13e44006
40060894
302c6057
36e461c3
40260215
4004303c
f32462d2
10944007
346f30ac
104c708c
3664306c
1110301c
0000311c
335c6c0c
04c307c4
40063664
0296552f
08040e56
0be5a0bc
00000804
fe961016
1110301c
0000311c
8c6c6c0c
6007710c
706c1b94
18546007
a6bc0fc3
40170bcd
640c306c
107423e4
069423e4
442c6057
30e402c3
001c0974
011c1150
28060000
26bc4006
029609d9
08040856
000620c3
31c32829
31a32849
31a32809
31a32869
31a32889
31a328a9
002662f2
00000804
0542041c
002602d2
00000804
ff967016
62c350c3
205c6364
8a6c0744
87d21fe6
015757ac
02c30037
466426c3
0e560196
00000804
50c33016
0744005c
04c382ac
17ac83d2
0c564664
00000804
305c20c3
335c0744
03c30844
0bac63d2
08043664
50c33016
0744005c
0d04405c
17ac83d2
0c564664
00000804
0be63cbc
00000804
1244305c
48bc63f2
08040be6
0be652bc
00000804
f7963016
41c350c3
21542007
20060fc3
a4bc4486
145c0bce
530c0e44
0d44345c
04156007
335c756c
80370e84
40b72077
345c60f7
61370dc4
0800343c
108c6177
70ac01b7
045c61f7
02370ee4
0784055c
82f21fc3
12bc14c3
09960bec
08040c56
0bd5ecbc
00000804
0bd804bc
00000804
0bd8c0bc
00000804
9ebc03ac
08040bc3
ff963016
42c3a117
406c4364
a03747d2
24c302c3
0bfaf2bc
a03700b3
28bc24c3
01960be6
08040c56
ff961016
803780d7
0be6acbc
08560196
00000804
fd96f016
62c370c3
20b71264
536453c3
0040253c
4c0f6217
1110301c
0000311c
335c6c0c
02c307a4
40c33664
27548007
4e097d6c
3f5c500d
702d0041
408c353c
41ac353c
60773364
00212f5c
6832504d
3f5c6037
706d0001
0040043c
16c3c6d2
b4bc25c3
00b30bcd
25c316c3
0bcea4bc
44d24257
0040343c
04c3680f
0f560396
00000804
fe961016
80378117
80778157
0be6cabc
08560296
00000804
0136f016
50c3fa96
72c320b7
832c83c3
22bc04c3
00070be6
80874a94
055c4854
52bc0784
0bd20be4
23c36097
07944027
65d2766c
0dc4335c
39546007
0380653c
10bc06c3
0fd20be6
00e04f3c
14c305c3
0be6a8bc
04c306f2
0be610bc
03d264c3
1140653c
01403f3c
60066037
05c36077
00412f5c
27c312c3
cabc38c3
40c30be6
15540007
60376157
16c305c3
888e201c
acbc34c3
50c30be6
1110301c
0000311c
335c6c0c
04c307c4
00533664
05c3bfe6
80760696
08040f56
00000804
00000804
00000804
00000804
00000804
08040006
00000804
09942127
111c301c
0000311c
335c6c0c
01930c84
0b3540a7
09b420a7
111c301c
0000311c
335c6c0c
36640ca4
00000804
00000804
00000804
00000804
00000804
00000804
00000804
00000804
00000804
00000804
00000804
00000804
00000804
00000804
00000804
00000804
0bc6a6bc
00000804
200c21c3
082f280f
442f200c
0804400f
bcbc002c
08040be7
602c200c
602c642f
60062c0f
602f600f
00000804
000620c3
32e4680c
00260294
00000804
1124305c
0c0c4c6c
08042664
305c1016
8dac1124
46640c0c
08040856
1344305c
6ad25fe6
111c301c
0000311c
335c6c0c
36640584
02c34006
00000804
0f36f016
a03c60c3
0ac32040
0be7d2bc
61940007
1104365c
5d946007
14c4365c
59946047
dabc06c3
01270be7
365c5494
60271524
331c0454
4d940080
1024565c
963c1410
b01c2800
b11c1110
08330000
0080753c
0fe4065c
400617c3
5ebc32c3
40c30be4
17c309c3
d2bc40c6
00070bcd
84d21e54
6007728c
05c31b54
0be7c8bc
111c301c
0000311c
335c6c0c
06c30564
265c17c3
36641224
1110301c
0000311c
335c6c0c
05c307c4
02b33664
06c387d2
243c17c3
e0bc0040
05c30be7
0be7c8bc
680c2bc3
07c4335c
366405c3
141058c3
bf945ae4
0f56f076
00000804
0336f016
71c360c3
43c382c3
1184105c
305c2fd2
6cd211e4
111c301c
0000311c
335c6c0c
005c0544
27c30fe4
80073664
465c3f54
963c1024
01332040
0080043c
40c617c3
0bcdd2bc
900c05d2
f79449e4
8bd20193
c8bc04c3
54c30be7
03e7831c
109110d4
01b354c3
babc0286
50c30bce
1e540007
17c30105
b4bc40c6
14910bcd
1024065c
748c0193
21c3208c
06d432e4
15c3002c
0be7bcbc
000c0113
f49409e4
15c3a4d2
0be7c4bc
f8bc06c3
c0760be7
08040f56
f8967016
51c340c3
63c302c3
145c4829
31c31344
309423e4
143c0045
d2bc2480
00070bcd
05c32994
2800143c
d2bc40c6
00070bcd
06c32154
13c37829
2fc32045
0be0c2bc
000720c3
045c1794
15c30fe4
5ebc32c3
07d20be4
6ed2628c
341c6117
6ad20001
15c304c3
03e8201c
341c6117
66bc0001
08960be8
08040e56
482c42ec
266402cc
00000804
30c31016
804c02ec
46640ecc
08040856
30c31016
808c02ec
46640ecc
08040856
40c31016
305c6006
628c0647
230c68d2
6c8c26d2
60063664
728f730f
08040856
600c24d2
03546027
62af6026
400f4026
305c6006
13c305a7
0cbc23c3
08040be9
40c31016
600c24d2
03546187
72af6026
500f4186
204604c3
04bc4026
04c30be9
400620a6
0be904bc
208604c3
04bc4026
60260be9
0607345c
08040856
40c31016
febc2026
00070be8
04c31154
febc20c6
0cd20be8
111c301c
0000311c
335c6c0c
04c30ce4
36642026
04c304b3
febc20c6
04d20be8
05c4345c
04c366d2
24bc2026
03130be9
05a4345c
0bf46647
12946667
345c6686
04c305a7
34bc2026
01530be9
111c301c
0000311c
335c6c0c
04c30d04
08563664
00000804
40c33016
6006a006
04c372af
0be952bc
63d272ac
ff13a026
0c5605c3
00000804
0804234f
0547105c
00000804
480c42ec
266402cc
00000804
02d230c3
03c3622c
00000804
602605d2
616660af
0804600f
40c31016
15540007
febc2006
00070be8
70ac1094
704c6ed2
60277fa5
724c0ab4
602663d2
04c3722f
40262006
0be904bc
08040856
05c7105c
00000804
101c07d2
111cf8e8
14bc0017
08040be9
0664305c
0014033c
00000804
40c31016
43a7402c
000c1494
f8f4101c
0017111c
0bcdd2bc
12ec0cf2
101c0ad2
111cf914
8ebc0017
04d20bce
00530026
08560006
00000804
40c31016
43a7402c
000c1494
f8f4101c
0017111c
0bcdd2bc
12ec0cf2
101c0ad2
111cf91c
8ebc0017
04d20bce
00530026
08560006
00000804
40c33016
06bc008c
a0060bcf
120cb08f
0bcf06bc
124cb20f
0bfb0cbc
04c3b24f
25c315c3
0be904bc
08040c56
000620c3
31c32829
31a32849
31a32809
31a32869
31a32889
31a328a9
002662f2
00000804
40a1041c
002602d2
00000804
0542041c
002602d2
00000804
0860041c
002602d2
00000804
0180041c
002602d2
00000804
1124305c
0c0c4c4c
08042664
1124305c
0c0c4c6c
08042664
1124305c
0c0c4c8c
08042664
fb963016
1124005c
8217a00c
82578037
82978077
82d780b7
831780f7
80cc8137
466405c3
0c560596
00000804
1124305c
0c0c4cec
08042664
1124305c
0c0c4d0c
08042664
ff963016
1124005c
8117a00c
812c8037
466405c3
0c560196
00000804
1124305c
0c0c4d4c
08042664
1124305c
0c0c4d6c
08042664
fe963016
1124005c
8157a00c
81978037
818c8077
466405c3
0c560296
00000804
005c1016
822c1124
4664000c
08040856
30c31016
1124005c
89d282ac
133c000c
233c0340
321c0240
466401e4
08040856
00000804
0f36f016
60c3ff96
92c381c3
e2d753c3
0184bf5c
0143af5c
32bc03c3
0ed20bea
2800463c
32bc04c3
08d20bea
14c306c3
0bea8abc
02740007
635754c3
12546007
111c301c
0000311c
43576c0c
435c4037
08c30444
27c319c3
46643bc3
00079fe6
bf5c1494
06c30007
2ac315c3
90bc37c3
40c30bea
111c301c
0000311c
335c6c0c
065c0424
36640fc4
1110301c
0000311c
335c6c0c
07c307c4
04c33664
f0760196
08040f56
01c330c3
335c2ad2
361c14e4
333c0001
7fe50b0d
03837f52
00000804
fb961016
1544305c
25946407
4007452c
654c2254
21946307
13c36809
433c6829
431c40ac
19b40fff
60376006
0020323c
20c66077
323c20b7
60f70080
41374206
201c2086
211cf924
34c30017
0bea6ebc
03740007
00530006
05961fe6
08040856
68bc2226
08040bea
00000804
40c31016
800701c3
00874354
00872f54
00270ab4
00071b54
00471454
00671f54
04331b94
2b5400e7
06b400e7
215400a7
129400c7
01070433
01272554
04b30d94
26544007
1447245c
323c0493
6c67fff0
245c1fb4
00061467
40070393
245c1954
ff531487
14c7245c
245cfef3
fe9314e7
1507245c
245cfe33
fdd31527
1547245c
245cfd73
fd131567
1587245c
1fe6fcb3
08040856
01e4021c
b4bc4106
08040bcd
40c3f016
52c371c3
24540007
1110601c
0000611c
335c780c
005c07c4
36641604
a8f2e2d2
345c6006
345c1607
03c31647
780c0253
07a4335c
366405c3
1607045c
17c309d2
b4bc25c3
545c0bcd
00061647
1fe60053
08040f56
40c3f016
52c371c3
24540007
1110601c
0000611c
335c780c
005c07c4
366415e4
a8f2e2d2
345c6006
345c15e7
03c31627
780c0253
07a4335c
366405c3
15e7045c
17c309d2
b4bc25c3
545c0bcd
00061627
1fe60053
08040f56
50c33016
000741c3
20073654
640c2454
1187305c
305c642c
644c11a7
11c7305c
305c646c
648c11e7
1207305c
305c64ac
24cc1227
021c2ad2
50ec0248
0bcdb4bc
355c70ec
00731347
1347105c
355c710c
02331367
1187155c
11a7155c
11c7155c
11e7155c
1207155c
1227155c
1347155c
1367155c
08040c56
40c37016
52c361c3
510f0cd2
0bcdb4bc
1767545c
2cc0043c
25c316c3
0bcdb4bc
08040e56
0136f016
40c3f796
72c381c3
636463c3
02003f3c
3f3c6037
607701c0
40062066
aabc6be6
50c30bea
a0071fe6
61d76454
14c4145c
20472177
201c0454
417700fe
00a11f5c
363c2c0d
273c0304
32a33005
61b73364
419761d7
41374832
00811f5c
61d72c2d
00c12f5c
345c4c4d
01d714c4
06946047
406d4006
4c8d61d7
006500f3
0030183c
b4bc4046
61d70bcd
0050033c
0050183c
b4bc4106
61d70bcd
135c2006
61d702ed
02f5135c
1524345c
643c01d7
42172800
4000331c
301c0e94
3f5c888e
a0770006
303c40b7
60f704d0
143c04c3
01b30d40
888e101c
00061f5c
40b7a077
04d0303c
04c360f7
0240143c
36c327c3
0bead4bc
80760996
08040f56
1f36f016
40c3f696
92c3a1c3
02a4bf5c
02e4cf5c
636463c3
02837f5c
81c32597
3f3c8364
60370240
02003f3c
20666077
383c4006
aabc05f0
50c30bea
a0071fe6
62176e54
14c4245c
404741b7
101c0454
21b700fe
00c12f5c
173c4c0d
363c2004
13a31085
621721f7
21772832
00a11f5c
62172c2d
00e12f5c
345c4c4d
021714c4
06946047
406d4006
4c8d6217
006500f3
0030193c
b4bc4046
62170bcd
0050033c
0050193c
b4bc4106
62170bcd
408c283c
1f5c4137
135c0081
621702ed
02c12f5c
02f5235c
68d23bc3
033c6217
1bc305f0
b4bc4597
345c0bcd
02171524
331c4257
0e944000
888e301c
00063f5c
40b7a077
04d0303c
04c360f7
03001c3c
101c0193
1f5c888e
a0770006
303c40b7
60f704d0
1cc304c3
3ac326c3
0bead4bc
f8760a96
08040f56
0336f016
70c3f396
82c351c3
605c2205
c1071504
4f3c1694
04c30140
b4bc4206
0f3c0bcd
153c0240
26c30280
0bcdb4bc
02c00f3c
0200153c
b4bc26c3
14c30bcd
14e4275c
746cd40c
95cc144c
0f944027
8f5c4037
00b70027
813720f7
16c307c3
6ebc4006
00070bea
02531515
4037542c
00278f5c
20f700b7
07c38137
201c16c3
211cf924
6ebc0017
00070bea
1fe60315
00060053
c0760d96
08040f56
40c37016
52c361c3
22540007
1110301c
0000311c
335c6c0c
005c07c4
366415a4
a8f2c2d2
345c6006
345c15a7
03c315c7
05c30213
0bfb26bc
15a7045c
16c309d2
b4bc25c3
545c0bcd
000615c7
1fe60053
08040e56
1f36f016
50c3f696
a2c3b1c3
c55783c3
02e4cf5c
a2dcc007
005c000c
50bc1524
40c30bea
32540007
155c0597
60801d64
0140033c
0bfb26bc
000740c3
000b72dc
459716c3
0bcdb4bc
111c301c
0000311c
335c6c0c
04c30e44
253c2597
36643400
26740007
6c006597
155c65b7
64c31d44
45972dd2
255c1100
b4bc1d64
65970bcd
1d64055c
65b76c00
259764c3
936491c3
02403f3c
3f3c6037
60770200
206605c3
393c4006
aabc05f0
70c30bea
301c0bf2
311c1110
6c0c0000
07c4335c
366404c3
62170eb3
14c4255c
404741f7
201c0454
41f700fe
00e10f5c
42170c0d
1085383c
420b033c
1f5c01b7
282d00c1
28c36217
41774372
00a10f5c
355c0c4d
021714c4
06946047
406d4006
4c8d6217
006500f3
00301a3c
b4bc4046
62170bcd
0050033c
00501a3c
b4bc4106
62170bcd
408c193c
2f5c2137
235c0081
621702ed
02c10f5c
02f5035c
033c6217
16c305f0
b4bc4597
301c0bcd
311c1110
6c0c0000
07c4335c
366404c3
033c6217
251700d0
b4bc4406
355c0bcd
02171524
331c4257
06944000
888e301c
00063f5c
101c00b3
1f5c888e
e0770006
303c40b7
60f704d0
1cc305c3
3bc328c3
0bead4bc
1fe60053
f8760a96
08040f56
50c3f016
42c371c3
1a540007
9ebc480c
00070be0
100f1574
15a4655c
c0076006
26bc1094
055c0bfb
0ad215a7
500c17c3
0bcdb4bc
355c700c
36c315c7
7fe60053
0f5603c3
00000804
10540007
1004105c
65ac28d2
2285610f
b4bc23c3
00d30bcd
610f6406
a4bc23c3
08040bce
0736f016
50c3fb96
83c3a1c3
01a49f5c
736472c3
04d0613c
00400f3c
420616c3
0bcdb4bc
0cc4355c
47546007
200606c3
a4bc4206
355c0bce
201c1524
211c111c
331c0000
08944000
c037680c
0444435c
1440053c
680c00f3
435cc037
053c0444
17c30640
39c328c3
0f3c4664
16c30040
d2bc4206
00070bcd
255c2094
32c31524
4000361c
0b0d333c
7f327fe5
0cc7355c
355c6026
231c0ca7
07944000
0a40053c
1140153c
00d34e06
0240053c
0640153c
b4bc4806
03f30bcd
0ca4355c
27546007
200606c3
a4bc4206
301c0bce
311c111c
6c0c0000
435cc037
053c0444
17c30240
39c328c3
0f3c4664
16c30040
d2bc4206
0df20bcd
1e40053c
00501a3c
b4bc4106
60260bcd
0f67355c
00530006
05961fe6
0f56e076
00000804
0336f016
50c3fd96
62c391c3
15e4305c
305c66f2
63f21604
0bea9ebc
0007180c
784c1994
23946007
15e4355c
355c65f2
60071604
382c1c54
40062037
786c4077
05c360b7
f92c101c
0017111c
600629c3
155c0a33
2bd215e4
455c582c
34c31624
209423e4
0bcdd2bc
1c940007
48c31850
25548007
1604755c
2154e007
1524055c
0bea50bc
111c301c
0000311c
255c6c0c
386c1644
435c2037
17c30504
466438c3
780c0ed2
4037582c
8077984c
20b7386c
101c05c3
111cf970
03730017
14c4355c
1c946027
4007584c
355c1954
60071604
355c1594
60071564
780c1154
8037982c
386c4077
05c320b7
f9ac101c
0017111c
64bc29c3
1fe60beb
055c02f3
50bc1524
00070bea
301c1054
311c111c
6c0c0000
0e24335c
19c305c3
366426c3
1fe630c3
02746007
03960006
0f56c076
00000804
ff967016
61c350c3
a4bc42c3
05c30bea
5cbc2126
80070bea
05c32154
406616c3
babc6026
055c0bea
20260fc4
0bfab2bc
1524055c
0bea4abc
055c06d2
20260fc4
0bfaa2bc
60376006
13c30026
ed3c201c
0017211c
3cbc35c3
255c0be5
45d21004
63d26a8c
6a8f6006
1524055c
0bea50bc
301c0bd2
311c111c
6c0c0000
0de4335c
200605c3
01963664
08040e56
40c3f016
000751c3
603c4c54
06c32800
b4bc40c6
043c0bcd
20061e40
a4bc4106
60060bce
0f67345c
345c6026
043c0f07
15c32180
d2bc40c6
0af20bcd
111c301c
0000311c
335c6c0c
04c30524
545c3664
a7d20c81
16c304c3
1cbc4026
04330bf0
111c701c
0000711c
335c7c0c
04c30dc4
00073664
045c1254
15c30fc4
0bfab2bc
16c304c3
1cbc4026
7c0c0bf0
0de4335c
15c304c3
00b33664
0ca7045c
0cc7045c
08040f56
41c37016
63c352c3
eebc01c3
41570be1
0ed2080f
e4bc04c3
61170be1
04c30c0f
0be1cebc
049450e4
65e40006
1fe60215
08040e56
0336f016
60c3ef96
72c391c3
8f3c43c3
08c30080
47862006
0bcea4bc
ffe0543c
35b4a407
243c47c3
323c011f
61770034
123c06c3
26bc088b
00f70beb
01800f3c
25c314c3
0bcdb4bc
265ca437
3f3c1504
60370100
00278f5c
12c306c3
35c325c3
0bf0b4bc
13940007
18c306c3
03d0293c
0bed70bc
0bf240c3
163c06c3
66172800
2004233c
0bf01cbc
005304c3
11961fe6
0f56c076
00000804
0136f016
50c3e596
43c3c857
8f3c4364
01c30080
28c312c3
0bde7cbc
3b740007
600761d7
34c33854
1000341c
33546007
433c6217
99cfffe0
1504255c
0080363c
c0776037
12c305c3
34c324c3
0bf0b4bc
000770c3
81d72094
32c35009
0003341c
7009786f
05c36232
0014133c
0beb26bc
6217182f
ffe0233c
0db44407
0100063c
0020143c
0bcdb4bc
18c305c3
0beb34bc
005307c3
1b961fe6
0f568076
00000804
0f36f016
a0c3f696
42c371c3
9f5cb3c3
6f5c02a4
44890283
446932c3
41ac823c
0dd139c3
32c344d7
68b443e4
c04754c3
80e70594
543c6335
3ac3ff80
1504235c
0080393c
9f5c6037
0ac30027
28c312c3
b4bc35c3
00070bf0
3b3c5194
29c3110b
c027686f
6f3c2994
06c30080
02d0173c
b4bc4206
0f3c0bcd
1a3c0180
42060340
0bcdb4bc
3ab48407
0100593c
173c05c3
24c305f0
0bcdb4bc
111c301c
0000311c
80376c0c
0484435c
240606c3
0100201c
466435c3
c0470333
343c2194
60070074
a4071d94
301c1bb4
311c111c
6c0c0000
0464435c
03400a3c
188c153c
05f0273c
0100393c
0af24664
1b3c0ac3
26bc098b
39c30beb
00060c2f
1fe60053
f0760a96
08040f56
0736f016
40c3ee96
83c352c3
0343af5c
0ce4305c
0001341c
5c546007
00c06f3c
200606c3
a4bc4786
04c30bce
0bea62bc
344990c3
342921c3
412c713c
02f1355c
355c13c3
233c02e9
345c40ac
604714c4
c0370994
153c04c3
37c305f0
0bf11abc
8f5c0173
af5c0007
c0b70026
15c304c3
6abc37c3
60c30bf1
210604c3
0bea5cbc
2894c007
1f3c04c3
253c00c0
70bc03d0
00070bed
04c31f94
2ac315c3
60bc37c3
00070bec
931c1774
09940009
a4bc04c3
04c30bea
5cbc19c3
01130bea
143c04c3
273c2800
1cbc2004
04c30bf0
0beac2bc
0f3c0173
200600c0
a4bc4786
04c30bce
68bc2026
12960bea
0f56e076
00000804
f996f016
61c350c3
21772006
005c21b7
002714e4
04bc5154
00070be2
055c4f54
eebc14e4
70c30be1
14e4055c
0be1cebc
055c40c3
e4bc14e4
355c0be1
163c14c4
604703d0
1f3c0394
355c0140
253c1524
331c2800
08944000
60376026
00b72077
0f40353c
602600f3
20776037
353c00b7
60f70440
05c38137
600617c3
0bea6ebc
1c740007
1364355c
16546007
111c401c
0000411c
0cec700c
400615c3
0be4e8bc
1364255c
6cec700c
20372006
23c302c3
3cbc35c3
00060be5
1fe60053
0f560796
00000804
0736f016
60c3e396
a2c371c3
20e6a364
0bea5cbc
9c49bc29
05f0073c
02f1275c
275c32c3
123c02e9
2f3c41ac
7cbc0100
00070bde
000963dc
422c853c
67d26257
341c38c3
60071000
0008c2dc
6bd26357
341c38c3
60071000
000842dc
63076397
000804dc
2800963c
19c306c3
01002f3c
0bef84bc
75740007
1bd0063c
00d0173c
d2bc4406
50c30bcd
6b940007
23c37c89
433c7c69
065c412c
cebc14e4
40e40be1
365c6094
331c1524
11944000
00068f5c
a0b7a077
0a40363c
06c360f7
27c319c3
debc3ac3
00070bec
02134c94
00068f5c
a0b7a077
0240363c
06c360f7
27c319c3
debc3ac3
00070bec
60263c74
0f07365c
0404383c
06c367d2
64bc17c3
00070bf2
383c3094
6cd22004
19c306c3
32c34026
0beababc
0fc4065c
b2bc2026
06c30bfa
5cbc2106
42570bea
8f5c4ad2
06c30007
629717c3
0bf0cebc
13740007
1f3c06c3
34bc0100
00070beb
62570c74
06c364d2
0beac2bc
0ce4365c
365c6072
00b30ce7
202606c3
0bea68bc
e0761d96
08040f56
0736f016
50c3ec96
82c3a1c3
2a544007
1004305c
c4dc6007
005c000e
5ebc0fe4
055c0be4
901c1007
00070001
000e14dc
08c31c33
42062085
0bcdd2bc
000740c3
05c31294
0beee6bc
111c301c
0000311c
335c6c0c
055c04e4
36640fc4
1767455c
98c31213
1524055c
0bea44bc
92dc0007
055c0008
00070fc4
000842dc
111c401c
0000411c
335c700c
15c304c4
36644406
0fc4255c
700c0bd2
04c4335c
15c302c3
36644206
63940007
700c03d3
00c06f3c
04c4335c
16c302c3
36644806
000740c3
000954dc
2cc0053c
02c01f3c
b4bc4406
44060bcd
1767255c
14c306c3
a4bc4806
10930bce
d50fc206
14c4355c
1f946047
1524455c
50bc04c3
00070bea
301c1894
311c111c
4c0c0000
0fe4155c
2700353c
355c6037
60771184
425c80b7
01c304a4
26c315c3
46643ac3
005360c3
383cc006
33c40b0d
f88c733c
1004455c
ebd28cf2
0fe4055c
28c31ac3
5ebc34c3
03d20be4
00f394c3
355cc6d2
63f21004
4294e007
1004355c
655c6ef2
01731007
1004355c
400665d2
1007255c
39c300f3
065365f2
400729c3
455c3154
04c31524
0bea44bc
2a540007
50bc04c3
20c30bea
24940007
04c03f3c
00776037
202605c3
aabc32c3
40c30bea
16540007
603764d7
153c05c3
201c2800
34c3888e
0bea90bc
1110301c
0000311c
335c6c0c
04c307c4
1fc63664
1fe601f3
000601b3
c4060173
901cefb3
155c0000
20071004
fff1d4dc
1496e693
0f56e076
00000804
0736f016
50c3fa96
82c391c3
305ca3c3
c60614e4
02946107
455cc806
04c31524
0bea50bc
0fd270c3
111c301c
0000311c
c0376c0c
0e64435c
19c305c3
3ac328c3
03b34664
56bc04c3
550c0bea
2800353c
353c6037
607719d0
00d0383c
af5c60b7
c1370067
05c30177
201c12c3
211cfa18
353c0017
e0bc2700
07c30be3
e0760696
08040f56
1f36f016
70c3e196
82c351c3
c364c3c3
0bea84bc
d2dc0007
07c3000b
5cbc20e6
4f3c0bea
04c30100
4c862006
0bcea4bc
14c4375c
12946047
05f0083c
325c28c3
63c302f1
02e9325c
123c23c3
24c3432c
0bde7cbc
93dc0007
07c30009
421715c3
0bf37ebc
52dc1fc7
00070009
0008e4dc
0f04375c
073c6bd2
240619d0
0bcecebc
34dc0007
075c0008
375c0f07
a73c1524
9f3c19d0
b73c0740
331c2800
3e944000
1140673c
200606c3
a4bc4e06
40060bce
0c27275c
111c301c
0000311c
335c6c0c
07c30404
26c318c3
573c3664
09c31740
410615c3
0bcdb4bc
17c0473c
14c305c3
b4bc4106
04c30bcd
410619c3
0bcdb4bc
375c6026
af5c0cc7
275c0007
407715a4
15c4375c
c0f760b7
1bc307c3
3cc328c3
0bede8bc
39940007
673c0613
07c30640
28c315c3
82bc36c3
573c0bf4
09c30940
410615c3
0bcdb4bc
09c0473c
14c305c3
b4bc4106
04c30bcd
410619c3
0bcdb4bc
275c4026
af5c0cc7
375c0007
607715a4
15c4275c
c0f740b7
1bc307c3
3cc328c3
0bede8bc
09740007
1bd0073c
00d0183c
b4bc4406
00b30bcd
202607c3
0bea68bc
f8761f96
08040f56
1f36f016
90c3ff96
62c3c1c3
200653c3
1c87105c
6c4741c3
000fd9dc
1110301c
0000311c
335c6c0c
05c307a4
b0c33664
00079fe6
000ef2dc
25c316c3
0bcdb4bc
0c493bc3
0c6910c3
233c30c3
0bc340ac
60676029
000d14dc
400ca23c
ffffa41c
408c323c
353ca3a3
a3e4ffc0
000c55dc
005ea31c
000c19dc
343c4bc3
331c021e
045400fe
84dc6047
29c3000b
0fc4025c
86bc2006
70490bfa
702903c3
402c733c
0074873c
0036383c
633c33c4
831cf88c
06540001
831cc5d2
04dc0002
29c3000a
1524525c
50bc05c3
05f20bea
56bc05c3
05d20bea
24dcc007
02530009
305c09c3
620714e4
831c0d94
0a540002
1504305c
42dc6207
373c0008
60070084
19c37f94
14e4315c
04946807
0002831c
09c37794
0f64305c
043c6ad2
193c0050
41061e40
0bcdd2bc
6af40007
341c37c3
60072080
373c6554
60078004
6a3c6194
a73c0040
2ac31004
c0374ad2
14c309c3
3bc328c3
0beef8bc
52940007
02f1345c
345c03c3
533c02e9
363c402c
53e4f9d0
19c347b4
14c4315c
19946047
341c37c3
60071000
301c1454
311c111c
6c0c0000
09c36fec
28c314c3
00073664
345c3194
03c302f1
02e9345c
402c533c
0084373c
14546007
0304373c
22946007
07d20ac3
14c309c3
c6bc28c3
03930bf2
1cc309c3
38c324c3
0bf4c4bc
37c302b3
2000341c
10946007
2ed21ac3
00068f5c
1cc309c3
35c324c3
0bf1ecbc
800600b3
9fe60093
80260053
1110301c
0000311c
335c6c0c
0bc307c4
04c33664
f8760196
08040f56
0be7f8bc
00000804
628c24d2
04546087
305c6026
40860607
6006428f
624f62ef
626f620f
612f614f
422f4026
00000804
628c24d2
04546107
305c6026
41060607
6026428f
0804630f
40c31016
63f2610c
6bf2618c
111c301c
0000311c
335c6c0c
04c30bc4
36642026
602773ac
60470454
00931194
6ed273cc
73cc0073
301c6bd2
311c111c
6c0c0000
0be4335c
200604c3
08563664
00000804
63ec24d2
045460c7
305c6026
40c60607
602643ef
0804620f
63ec24d2
045460e7
305c6026
40e60607
602643ef
0804626f
63ec24d2
04546047
305c6026
40460607
600643ef
4026622f
0667205c
00000804
40c33016
0864305c
0cccad0c
201c2046
211cfa30
60060017
345c5664
602504e4
04e7345c
04a4345c
345c6025
0c5604a7
00000804
0864005c
64d2624c
2026000c
08043664
40c31016
628c24d2
04546127
345c6026
41260607
6026528f
04c371af
0bf72cbc
532f4046
08040856
40c31016
628c24d2
045460a7
345c6026
40a60607
6026528f
04c371af
0bf72cbc
245c4026
08560887
00000804
0864005c
64d2624c
2006000c
08043664
40c31016
628c24d2
04546047
345c6026
40460607
04c3528f
0bf712bc
72cf6026
51af4006
5ebc04c3
08560bf7
00000804
40c31016
628c24d2
04546147
345c6026
41460607
6006528f
04c371af
0bf75ebc
532f4026
12bc04c3
08560bf7
00000804
40c31016
628c24d2
04546027
345c6026
40260607
6006528f
72ef732f
71af72cf
5ebc04c3
40260bf7
600651ef
08c7345c
08e7345c
0856702f
00000804
305c06d2
602504a4
04a7305c
00000804
2d540007
1d542087
09b42087
12542027
20472fd2
20671154
02132294
175420c7
121420c7
155420e7
19942107
00ec02b3
030c02f3
00ac02b3
005c0273
02130444
0404005c
005c01b3
01530424
0113018c
06e4005c
005c00b3
00530704
08040006
2c540007
1d542087
09b42087
12542027
20472fd2
20671154
02132194
175420c7
121420c7
155420e7
18942107
40ef02b3
430f02b3
40af0273
205c0233
01d30447
0407205c
205c0173
01130427
00d3418f
06e7205c
205c0073
08040707
23f204d2
0053006c
08040006
0007fe96
20ec1054
2df22077
00213f5c
60ac23c3
402662f2
0016323c
0f5c6037
00530001
02960006
00000804
40c33016
000752c3
105c2154
40070647
680c1d54
07c7305c
305c682c
684c07e7
0807305c
305c686c
005c0827
0ed20624
a0bc284c
045c0be9
346c0624
0be9a2bc
0624045c
d2bc348c
0c560be9
00000804
ff963016
a08c40c3
1594a007
608f6026
f584001c
0017011c
24c315c3
0be4e8bc
00268037
201c15c3
211cf584
35c30017
0be53cbc
0c560196
00000804
25f206d2
43d2406f
0bf85ebc
00000804
40c31016
628c24d2
045460e7
345c6026
40e60607
734c528f
04c3702f
0bf85ebc
51af4006
5ebc04c3
60460bf7
0887345c
08040856
40c31016
4bd242ac
69f262cc
67f2610c
65d2618c
66bc2026
18530bf7
23f2316c
65f2732c
63f2710c
64f2718c
202604c3
204705f3
732c0994
0f546047
202604c3
0bf734bc
202715b3
732c0894
05546027
7ebc04c3
14930bf7
6087728c
60874c54
604709b4
60471054
602716b4
000994dc
60e70d93
61077454
0008e2dc
04dc60a7
0f930009
c4dc4007
04c30008
96bc12c3
10d30bf7
4007504c
72ec1694
01c3338c
0c3430e4
111c301c
0000311c
335c6c0c
04c30d24
366412c3
71cc0e73
04c364d2
065312c3
63f270ec
24d230ac
200604c3
70cc0cb3
600704c3
40075794
72ec6194
01c3338c
5c1430e4
600771cc
04c35994
04b312c3
600770ec
71cc1154
345c6ff2
6cd207c4
07e4345c
202669f2
045c31cf
60ec0864
000c63d2
70ec3664
71cc68d2
04c366d2
48bc2006
07530bf7
65f270ac
68d2712c
66f271cc
200604c3
0bf884bc
726c05f3
2c546007
111c301c
0000311c
335c6c0c
04c30d24
f5d32006
2af2302c
111c301c
0000311c
335c6c0c
04c30d24
70ccf473
14546007
70cc00b3
71cc68d2
04c366d2
b6bc2006
01530bf6
04c331cc
efd327f2
24f2330c
a2bc04c3
08560bf6
00000804
40c31016
63ec24d2
04546107
345c6026
41060607
602653ef
724f714f
0624045c
0be9acbc
400604d2
0727245c
08040856
40c33016
0684005c
0bfb0cbc
545ca006
045c0687
06bc06c4
545c0bcf
045c06c7
1cbc0624
0c560bea
00000804
40c31016
63ec24d2
04546027
345c6026
40260607
04c353ef
0bf988bc
71ef6006
0856700f
00000804
20c31016
63f2610c
26d221ec
202602c3
0bf99ebc
63ec0ed3
59546087
08b46087
36546047
0db46047
6b946027
60c709b3
60c74b54
60e72514
61074754
08936294
0444405c
301c89d2
311c111c
6c0c0000
0d44335c
105c0193
2bd20404
111c301c
0000311c
335c6c0c
14c30d64
09333664
600760ac
60ec3994
43546007
301c0453
311c111c
6c0c0000
0d64335c
60acfe13
622c64d2
28946007
6dd268cc
6bd26a2c
111c301c
0000311c
335c6c0c
02c30d84
fbb32006
600768ec
6a2c2454
21546007
200602c3
02bc0393
03730bf7
69d260cc
111c301c
0000311c
335c6c0c
f8f30d84
85d280ac
eabc13c3
01730bf6
24f2200c
0bf6f6bc
60ec00d3
14c364d2
0bf970bc
08040856
ff963016
800650c3
355c6006
05c30607
0bf89ebc
c2bc05c3
05c30bf6
0bf9b2bc
0624055c
0be990bc
602604d2
0607355c
0604355c
802564d2
e7948c87
0604355c
13546007
f57c001c
0017011c
25c32006
0be4e8bc
0006a037
201c10c3
211cf57c
30c30017
0be53cbc
0864355c
60076c4c
155c1754
20070884
20271354
055c0854
debc0624
20460be9
10c302f2
355c6006
355c0887
8c4c0864
4c6c05c3
01964664
08040c56
40c33016
09d251c3
0624005c
0be9b8bc
04c3a4f2
0bfa34bc
08040c56
216f04d2
0bfa34bc
00000804
20af06d2
0707105c
0bfa34bc
00000804
40c31016
20ef0cd2
06e7105c
005c25d2
b2bc0624
04c30be9
0bfa34bc
08040856
21cf04d2
0bfa34bc
00000804
218f04d2
0bfa34bc
00000804
34bc01c3
08040bfa
ff963016
41c350c3
63d2640c
640f7fe5
63d2702c
702f7fe5
63d2704c
704f7fe5
63d2706c
706f7fe5
500c702c
504c32a3
506c32a3
6cd232a3
00268037
201c2006
211cf584
35c30017
0be53cbc
708f0053
34bc04c3
01960bfa
08040c56
08040006
08040006
08040006
00000804
08041fe6
00000804
c4bc1016
40c30a80
301c09f2
311c0b84
6c0c0000
220c001c
04c33664
08040856
18540007
8000101c
fbc1111c
201c6080
211cafff
12c30000
0ab431e4
0b84301c
0000311c
001c6c0c
366422a8
5cbc0073
08040a7f
40061016
0ff402e4
0a7e8abc
20c340c3
301c0af2
311c0b84
6c0c0000
2222001c
24c33664
085602c3
00000804
0136f016
fdecf21c
51c340c3
83c362c3
0005831c
0fc321b4
25c314c3
26bc36c3
00070b1d
40c31994
0fc301d3
11643f5c
4a1d133c
11843f5c
4a1d233c
0b1d14bc
80250bf2
f21448e4
1f5c0fc3
04bc11a4
30c30b1d
1fe662d2
0214f21c
0f568076
00000804
fd967016
51c340c3
603762c3
607761d7
60b76217
14c30026
36c325c3
0bfb3cbc
0e560396
00000804
40f7fc96
3f3c60b7
60370080
60776157
3f3c4026
6ebc00c0
04960bfb
00000804
0bfb0cbc
00000804
0bfb0cbc
00000804
12c331c3
52bc23c3
08040a9c
ff967016
61c350c3
0130001c
0bfb26bc
20c340c3
20260fd2
15c32037
600626c3
0b1e8cbc
000724c3
04c30515
0bfb0cbc
02c34006
0e560196
00000804
ff967016
61c350c3
0130001c
0bfb26bc
20c340c3
20060fd2
15c32037
600626c3
0b1e8cbc
000724c3
04c30515
0bfb0cbc
02c34006
0e560196
00000804
12c331c3
3ebc23c3
08040aa1
01f25000
00000001
00307061
6d206f6e
68637461
206e6920
6e616373
00000000
45524944
002d5443
5f617077
5f737362
6f6d6572
6f5f6576
7365646c
00000074
5f617077
5f737362
6f6d6572
6f5f6576
7365646c
6e755f74
776f6e6b
0000006e
ffffffff
0000ffff
5f617077
70707573
6163696c
7620746e
0a302e32
79706f43
68676972
63282074
30322029
322d3330
2c323130
756f4a20
4d20696e
6e696c61
3c206e65
3177406a
3e69662e
646e6120
6e6f6320
62697274
726f7475
00000073
73696854
666f7320
72617774
616d2065
65622079
73696420
62697274
64657475
646e7520
74207265
74206568
736d7265
20666f20
20656874
20445342
6563696c
2e65736e
6565530a
41455220
20454d44
20726f66
65726f6d
74656420
736c6961
00000a2e
61766e69
6164696c
00006574
2d414657
706d6953
6f43656c
6769666e
726e452d
656c6c6f
2d312d65
00000030
3d6e6970
00000000
3d636270
00000031
ffffffff
0000ffff
69204549
2f33206e
736d2034
6f642067
6e207365
6d20746f
68637461
74697720
45492068
206e6920
63616542
502f6e6f
65626f72
70736552
6f6e2820
3f454920
00000029
69204549
2f33206e
736d2034
6f642067
6e207365
6d20746f
68637461
74697720
45492068
206e6920
63616542
502f6e6f
65626f72
70736552
00000000
73736f50
656c6269
776f6420
6172676e
61206564
63617474
6564206b
74636574
2d206465
4e535220
73617720
616e6520
64656c62
646e6120
4e535220
20454920
20736177
6d206e69
33206773
202c342f
20747562
20746f6e
42206e69
6f636165
72502f6e
5265626f
00707365
72696150
65736977
79656b20
70786520
69736e61
00006e6f
00000000
00000004
fc967016
20372066
f88c603c
404604f2
03734037
cbd240c3
600640c4
cf00311c
111c2006
21c38000
145402e4
a0b7a3c6
04c380f7
0a9428bc
00071fe5
343c06f4
60f7000d
60b77420
0fc3c077
0bfd4abc
03c330c3
0e560496
00000804
406c3016
600ca02c
03b46027
09335472
46546087
04946047
12c34006
12c30893
41544007
1047004c
70462715
00066c20
0cd46327
308d123c
343c8026
033c300d
0283fff0
04c302d2
303c01a3
680707f4
303c0694
64d20804
00530805
200607e5
ffff301c
3fff311c
02e423c3
20260235
388c203c
0fe70313
103c13d4
323c07f0
680707f4
323c0694
64d20804
00534805
400747e5
41320315
47322025
40060093
00ff101c
ffff001c
007f011c
253c2083
313cf92c
033c0ff4
0c56b92c
00000804
140460c3
00000804
08041fe6
14b8301c
0000311c
4c0f4186
08041fe6
14b8301c
0000311c
4c0f4166
08041fe6
2000301c
0006642f
00000804
08040026
08040026
14b8301c
0000311c
4c0f42c6
08041fe6
14b8301c
0000311c
4c0f43e6
08041fe6
08040006
08041fe6
08040006
20c31016
14b4001c
0000011c
6007600c
301c1954
311c14b0
000c0000
2c0c4100
24e441c3
301c07b4
311c14b4
4c0f0000
301c0313
311c14b8
21860000
1fe62c0f
101c0213
111c0004
200f0018
14b0301c
0000311c
0004401c
0018411c
fbd38c0f
08040856
2000301c
0006642f
00000804
08041fe6
14b8301c
0000311c
4c0f4046
08041fe6
14b8301c
0000311c
4c0f4146
08041fe6
08040006
68d230c3
14b8301c
0000311c
4c0f4b06
08041fe6
14b8301c
0000311c
4c0f4b06
08041fe6
50c33016
42c301c3
2b544007
35a331c3
0003341c
fff0123c
28946007
806715c3
540c2235
53c3600c
185425e4
501c0393
511cfeff
6a80fefe
328322e3
8080201c
8080211c
6df23283
00852085
1c358067
a00c440c
23e435c3
9f850694
e8948007
03130006
143c51c3
7408fff0
23e44008
37d20e94
353c56d2
203c008e
23e4008e
3fe50694
51c3fef3
ee948007
60095409
0c5609a0
00000804
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
c8134fb1
1ee2f1fe
