10fc301c
0000311c
00064c0c
6c6c704c
029434e4
696c0026
506c3664
084f104c
4c6f704c
342c702c
742f6c80
301c9580
311c10fc
4c0c0000
702c0006
021530e4
696c0026
142c3664
373c100f
62d24004
0f56f324
00000804
60c3f016
13bc401c
0000411c
500f4006
904f502f
31c3906f
32835f86
ff80733c
10fc501c
0000511c
27e3740c
023c6d6c
3664f88c
780f6006
03c3b40c
6c4c706c
31e414c3
00260294
3664756c
10fc301c
0000311c
00064c0c
13bc301c
0000311c
6c6c6c4c
13bc401c
0000411c
31e414c3
00260294
3664696c
13bc301c
0000311c
4c6c784f
cc6f586f
cc4f786c
9b80f82f
301cf00f
311c10fc
6c0c0000
00266d6c
60063664
8000311c
0f56702f
00000804
61c3f016
201c52c3
211c13bc
884c0000
13b4201c
0000211c
2c0f280c
13b8301c
0000311c
41572c0c
301c280f
311c13ac
4c0c0000
6006400f
3fe6780f
701c340f
711c10fc
02930000
00065c0c
30e4702c
002602f4
3664696c
502c780c
780f6d00
340c702c
32e421c3
740f02f4
301c904c
311c13bc
13c30000
e79441e4
08040f56
60c3f016
01c351c3
0a7e8abc
000770c3
c0071f54
365c1d54
33c4ffe4
ff80433c
10fc301c
0000311c
343c4c0c
6e20f90c
033c496c
2664f88c
45e424c3
25c302f4
16c307c3
08cbb0bc
5cbc06c3
07c30a7f
08040f56
60c37016
0a7e8abc
000740c3
305c1b54
33c4ffe4
ff80533c
305c65f2
533cffa4
301cff40
311c10fc
6c0c0000
56e40006
00260274
36646d6c
200604c3
b0bc25c3
04c30891
08040e56
2049fe96
20072077
60691294
0f946807
00213f5c
608923c3
0096331c
40260254
0016123c
0f5c2037
00530001
02960006
00000804
20c33016
426441c3
692c0b85
01732180
35c3ac09
41806045
09b421e4
34e46009
02c30754
0010303c
f31431e4
0c560006
00000804
11643016
436442c3
63d2632c
329460a7
0764305c
40474c4c
20072d94
ae242674
002cf524
0101305c
301c6df2
311c1110
6c0c0000
0404335c
101c04c3
36644321
305c01f3
6cd20101
1110301c
0000311c
335c6c0c
04c30424
4321101c
353c3664
68d24004
00d3f324
6d4c62cc
27e602c3
0c563664
00000804
3f36f016
82c341c3
40102330
a2d08030
0293b15c
62ac0ac3
04c4735c
0001931c
500b0994
321c32c3
501c00ff
3583ff00
931c0133
07940002
30c3100b
3f866065
700e3183
500b904f
336432c3
0200331c
201c0335
50ce0200
b300d02b
60077489
d5801c54
20061b80
00735780
600d68a2
1fe53fe5
60076780
56c3fa15
f02bd889
702e7b80
233c740c
1489600b
323c4820
740f601b
348d2006
0283345c
233c540c
540f231b
0283345c
719460a7
60277449
7cc36e54
035c7e0c
00070669
1ac36894
635c66ac
570004c4
a7c3e909
373ce929
0889452c
08a910c3
40ac603c
6ca034eb
736473c3
1110301c
0000311c
2c0c6c0c
a0c30849
303c0869
333c452c
442c03c7
6e696d00
059460c7
61cc0dc3
366404c3
233c740c
7f00fff4
395423e4
1954e6c7
35b4c247
0001b31c
301c0935
311c0b84
6c0c0000
4201001c
100b3664
7dc57800
30cb700e
7dc57880
163c70ce
0313fee0
1db4c0c7
0001b31c
301c0935
311c0b84
6c0c0000
4202001c
f00b3664
7f457b80
10cb700e
7f457800
163c70ce
740cffa0
600b233c
323c4500
740f601b
0b0d393c
233c7fe5
393cf88c
333c0026
7fe50b0d
f88c533c
a7f248f2
0006931c
25c30454
085315c3
38c3d04c
0006cc0f
0006931c
20860554
204e08c3
44f20026
0006931c
702b0a94
d80c68c3
78c36f00
0f9d373c
02734006
31c3302b
fffc341c
480c28c3
68c36d00
0f9d363c
37c3f02b
0003341c
7f3233c4
080c233c
303c2364
68c3180c
f0cb3980
7f20d02b
644e6980
0010103c
37c3f00b
102b6085
69806c20
323c700e
702e0040
323c4026
63120010
313c1180
48c3180c
01337180
cc0fc00c
ec4ee04b
20254025
61050105
f7142be4
313cabd2
7f05180c
418008c3
34c3884b
bf866065
931c0213
0f940001
7ca079c3
1b0c333c
418008c3
34c3884b
00ff321c
ff00501c
684e3583
180c313c
198068c3
0f56fc76
00000804
3f36f016
301cff96
311c0bb4
8c300000
0804635c
22100cc3
701ca006
711c1110
b3c30000
0ef0d01c
0000d11c
78bc0126
982c08cc
79548007
145c2006
109004a7
62f2780c
7fe51004
782c780f
782f6c0c
784f62f2
82bc0126
345c08cc
608701d1
39c31d94
0681335c
7c0c69f2
044918c3
36646fcc
516450c3
7c0ca9f2
04c36fec
03643664
0007a006
2dc3d294
1bc3680c
143c040c
36640040
60a7f953
5c0c4394
6d2968cc
0d946027
21c909c3
21e981c3
303c01c3
65f2442c
0444325c
366404c3
01c3a45c
66ec1bc3
508c0f10
335c39c3
00260669
10946007
662c1cc3
70126d69
011c0006
30830004
28496dd2
20272037
0f5c0994
084d0001
6f6c7c0c
366404c3
7c0c00f3
04c36dcc
50c33664
001c5164
011c0bb4
15c30000
28a42ac3
0a8146bc
1004f0d3
f0731004
82bc0126
019608cc
0f56fc76
00000804
fe96f016
51c360c3
802ce32c
6cec616c
36640006
226420c3
0301345c
13546007
1154e007
0f54e087
cccc101c
0000111c
0407155c
00d0301c
2100311c
33646c0b
0427355c
2954e087
0101345c
05356027
01d1355c
0b5460a7
01d1355c
1d946087
6c2c780c
6c2b6c2c
17b460c7
4c6c780c
03c34a4c
0040153c
e4d22664
74dce0a7
365c0008
0c4c0764
14dc0047
7acc0008
27e66d4c
0f733664
0101345c
345c6dd2
133c0101
20370010
00013f5c
0f5c6077
045c0021
40070105
580c1154
6e4c686c
153c02c3
36640040
8d6c7acc
00a5001c
49e62006
46646006
355c0b53
60a701d1
720c3394
0669035c
2e540007
04a7255c
1110301c
0000311c
68cc4c0c
60276d29
720c0c94
10c30dc9
303c0de9
65f240ac
0444325c
366405c3
378b7aec
65204f0c
436443c3
0026748c
301c0c4d
311c1110
6c0c0000
05c36f6c
06c33664
24c32006
0a8146bc
01260493
08cc78bc
0804365c
40254c0c
265c4c0f
684c0804
a82f63f2
ac0f0053
0804365c
365cac4f
6c4c0804
2c0f2006
82bc0126
008608cc
301c2066
311c0fe4
4d0c0000
08c8d4bc
0f560296
00000804
3f36f016
70c3d396
62b7a1c3
b364b2c3
21c32289
313c22a9
42c9412c
81ac323c
043c82e9
175cc1ac
21c305e9
05f1175c
412c313c
05f9275c
81ac323c
0601475c
c1ac143c
301c22f7
311c1110
4c0c0000
0764125c
600623b7
058d3f5c
4f5c81e6
35860595
059d1f5c
05753f5c
3f5c6a06
4bc3057d
82dc8007
00070028
002852dc
1f5c2886
6926053d
05453f5c
4f5c8a46
28a6054d
05551f5c
3f5c6866
8a86055d
05654f5c
1f5c25a6
7e46056d
05853f5c
00a01a3c
da3c2337
4ac30100
31c33009
00f0341c
0080331c
331c1854
08b40080
b2dc6807
6a070024
002594dc
331c01d3
72dc00c0
331c0024
82dc00d0
331c0022
c4dc00a0
48330024
0161275c
275c42c3
323c0169
475c422c
343c0171
075c81ac
903c0179
b31cc1ac
69dc0024
3b3c0023
c3c3fdc0
9e49c364
9e6904c3
402c343c
0b946027
02600a3c
0a701f3c
eabc40e6
000708cb
002234dc
21c33dc9
313c3de9
6007412c
0a3c1154
173c0260
375c0360
43c302b9
02c1375c
422c233c
0bcdd2bc
c4dc0007
a0060020
02608a3c
800749c3
40933294
100c653c
600c09c3
5a1d033c
2cbc2006
04f20a81
40c30377
403c00b3
00290020
19c30377
6f01640c
0530033c
40c61dc3
08cbeabc
11940007
18c304c3
01a13f5c
2abc23c3
01640892
49c308f2
cf01700c
d4dcc007
0153000b
0010353c
536453c3
202c09c3
52e421c3
39c3cc14
501c2c2c
511c1110
21470000
000849dc
435c740c
29c30864
4086080c
46646397
49c36026
6e20902c
400c09c3
130c333c
6cec6981
21c32e17
127432e4
05b9475c
475c04c3
343c05c1
6007402c
0dc34054
0300173c
eabc40c6
000708cb
075c3894
10c305b9
05c1075c
40ac303c
22546007
19c36026
6ca0242c
500c49c3
130c333c
033c6981
173c0530
40c60300
08cbeabc
10940007
133c702c
2277ffe0
533c700c
74ec1a1d
01216f5c
42c34e17
11f434e4
09c32eb3
313c202c
400c100c
a9817f85
fff0313c
6f5c6237
00730101
65c3a006
1110801c
0000811c
700c48c3
0784335c
05c00c3c
40c33664
82dc0007
acd20015
600c08c3
07c4335c
366405c3
640c19c3
6b9d433c
28c308f3
335c680c
366407c4
28b305c3
335c740c
0c3c0784
366405c0
000760c3
0013b2dc
49c3540c
6025702c
07e4225c
133c100c
2664100c
08f240c3
335c740c
06c307c4
04c33664
09c32513
643c602c
602c3b9d
602f6025
0373800f
1110801c
0000811c
640c18c3
0784335c
05c00c3c
40c33664
02dc0007
28c30011
335c680c
06c307c4
09c33664
433c600c
64c35b9d
25f22297
00ad001c
0a7762bc
0530063c
40c61dc3
08cbb0bc
0140063c
01801a3c
b0bc4106
429708cb
3f5c582f
365c0721
0dc3016d
0300173c
eabc40c6
0cf208cb
04c48e17
0f5c01f7
075c00e1
165c0a15
175c0169
2ac30a0d
588e4a0b
722b4ac3
993178ae
18ef0e17
41b720c4
00c14f5c
017d465c
341c23c3
68d20001
0024323c
002665f2
0185065c
20060093
0185165c
32c358ab
0010341c
65d26177
465c8066
00b30175
00a10f5c
0175065c
05c0063c
02401a3c
b0bc2cc3
06c308cb
2cbc2006
0ed20a81
463ca029
04c30310
9cbc2446
04c308cb
02601a3c
b0bc25c3
848608cb
0ae08f3c
a6001ac3
6622f429
00dd331c
05c32c94
0a8112bc
602605d2
0165365c
343c0493
1ac30020
18c30580
eabc4066
000708cb
54a91a94
40274137
0f5c1694
065c0081
243c0175
74cb00e0
49806212
65621ac3
65806212
41176d00
60276d22
20860494
0175165c
0020373c
43c37180
4be44364
06c3c814
2cbc2606
40c30a81
14540007
1f3c0085
40660b10
08cbeabc
60460df2
0175365c
6212708b
6de97180
04946027
065c00a6
22d70175
01c327d2
23170305
eabc40c6
301c08cb
311c1110
6c0c0000
0864435c
0c0c39c3
40862c2c
46646397
b31c0533
24350019
27091ac3
00051f5c
01903a3c
3b3c6077
60b7fe70
60f76297
0824425c
00401a3c
3dc34317
02534664
0018b31c
01930fb4
0844325c
009321a6
0844325c
2f3c2026
366403c0
1fc60073
00060053
fc762d96
08040f56
301cf016
311c1114
6c0c0000
ee24ac6c
4004673c
0046f524
08cc78bc
6af2746c
82bc0046
373c08cc
60074004
f3241954
948c02f3
004688f2
08cc82bc
1054c007
01d3f324
746f7fe5
748f702c
82bc0046
c2d208cc
04c3f324
0bc2f8bc
0f56fb93
00000804
50c37016
28540007
f524ce24
1114301c
0000311c
8c6c6c0c
600f6006
78bc0026
702c08cc
704c64d2
0053ac0f
b04fb02f
6025700c
0026700f
08cc82bc
20460066
0fe4301c
0000311c
d4bc4d0c
363c08c8
62d24004
0e56f324
00000804
301c3016
311c0bb4
8c2c0000
1110501c
0000511c
6d6c740c
720c3664
07c9135c
720c2bf2
12c34dc9
323c4de9
64f240ac
6d2c740c
0c563664
00000804
301c7016
311c0bb4
ac2c0000
1110301c
0000311c
c46c2c0c
4c6c766c
1a944007
86a0001c
0001011c
301c254c
311c0b54
5abc0000
201c0874
211c10f0
680c0000
680f6025
10ee201c
0000211c
6025680c
401c680f
411c10f0
700c0000
22356127
10f4101c
0000111c
700c040c
141d4146
6c003320
700c640f
3320341d
762c700f
78126e09
211c4006
32831000
560c6bd2
1110301c
0000311c
6d8c6c0c
1550023c
790c3664
786c6df2
782c64f2
08f46007
1110301c
0000311c
6dac6c0c
0e563664
00000804
41c33016
642f6006
53c36e24
f5245364
78bc0e26
201c08cc
211c0ef4
680c0000
680f6025
63f2684c
0053882f
301c8c2f
311c0ef4
8c4f0000
702f6006
82bc0e26
301c08cc
311c0bb4
6c4c0000
2c0c0046
0fe4301c
0000311c
d4bc4d0c
353c08c8
62d24004
0006f324
08040c56
1150001c
0000011c
40062406
09d926bc
00000804
1150001c
0000011c
404637e6
09d926bc
0be5e4bc
00000804
1150001c
0000011c
40463be6
09d926bc
0a82d4bc
00000804
1150001c
0000011c
40463de6
09d926bc
0a8704bc
00000804
60b7fd96
602764d2
02f32794
23c368a9
40775fc5
00213f5c
04356027
602761e9
40260694
716644cd
02d3650d
04cd0026
00412f5c
0213450d
03c368a9
00371fe5
00013f5c
08b46047
00413f5c
680c64cd
01e1035c
0396050d
00000804
3f36f016
70c3fd96
82c3c1c3
901cc00c
911c1114
19c30000
ac50640c
535c888c
14c30544
602626c3
2dc35664
b4c36aac
0484135c
700cb184
323c43c6
4086601b
231b323c
4006700f
6306504d
19c370ad
a35c640c
7c0c0564
586bac0c
0010323c
cf5c786e
2f5c0007
201c0026
2f5c013a
0bc30046
2cc33606
0010353c
3bc3a664
125c5c0c
133c0453
40260c6e
20064c2e
3dc32c4e
700c4eac
0fff341c
0484125c
33646c80
68ce28c3
19c36b8e
6d2c640c
366408c3
fc760396
08040f56
62c3f016
526451c3
436443c3
01734006
20291900
35e46009
313c0954
69800020
236423c3
f51424e4
0f560006
00000804
fe963016
31c320c3
45b9415c
08b8101c
20060c80
01b32264
013f303c
049432e4
20772026
513c0153
a0370010
00011f5c
f31414e4
a077a006
00211f5c
029601c3
08040c56
c00cf016
442bb80c
2c896500
420521c3
5c09ed00
341c32c3
43c30001
17946007
07c301b3
0010153c
eabc40c6
0ad208cb
0010343c
436443c3
365cab85
34e403a3
365cf1b4
04c303a3
029434e4
0f561fe6
00000804
0736f016
50c3fe96
42c381c3
af5c93c3
642b0143
ec80244c
61ccc00c
0001341c
78a96ad2
07946027
0823105c
602531c3
0826305c
1114301c
0000311c
6c0c6c0c
335c6c0c
620703e3
78a91894
03546027
13946067
00a0043c
6ba0163c
eabc40c6
0bf208cb
0040043c
0150153c
eabc40c6
03f208cb
4526065c
1114301c
0000311c
680c4c0c
335c6c0c
610703e3
62071254
78a95d94
165c65d2
2bf24543
325c0af3
1de90584
366416c3
326430c3
4e546007
602778a9
60670654
80060454
1b946007
1114301c
0000311c
5de96c0c
00052f5c
115c18c3
1f5c0681
8f8c0025
193c05c3
40060100
ff003a3c
40c34664
00264164
2d748007
62d72026
55462c0e
7de95c4d
701c7d0d
711c1114
7c0c0000
08c36dcc
80473664
55091b94
742c4dd2
03e3335c
08946207
566d5629
335c7c0c
05c30504
301c3664
311c1114
6c0c0000
8e4cc037
20060266
600621c3
00064664
e0760296
08040f56
0f36f016
fdf0f21c
61c390c3
844c642b
a0064e00
10765f5c
0021a25c
b33c680c
8849fff4
01003a3c
838482c3
480928c3
301c40b7
311c1178
5f5c0000
ac0d0041
0b548047
1114301c
0000311c
335c6c0c
2f3c0464
0db300e0
43c36097
0080431c
53c31154
2a0713c3
23c30d54
44076bd2
a6070954
a0060754
00e07f3c
420723c3
48c32294
b8cb7320
53c375a0
365c5364
78c30293
17356027
00e04f3c
18c304c3
b0bc25c3
594b08cb
74c37500
0200331c
12800ad4
b0bc388c
594b08cb
53c37500
74c35364
1178301c
0000311c
6a076c09
201c1854
211c1114
331c0000
23940080
fe803b3c
5f5c480c
3aa40006
00263f5c
09c38a2c
28c316c3
466437c3
1c940007
1114301c
0000311c
5f5c4c0c
3f3c0006
607720e0
04a4425c
16c309c3
37c328c3
01534664
335c680c
09c30464
27c316c3
01643664
4f5c02f3
00061073
12948007
1114301c
0000311c
6c4c6c0c
235c6c6c
301c05a4
311c0bb4
0c0c0000
266416c3
f21c04c3
f0760210
08040f56
40c3f016
7f5c53c3
6f5c00c3
200d00e3
602d6006
12c30085
b0bc40c6
043c08cb
15c300a0
b0bc40c6
043c08cb
21570100
b0bc40c6
d02e08cb
200c373c
0f56716e
00000804
0136f016
51c370c3
301c5264
311c1114
6c0c0000
301c0c50
311c1110
6c0c0000
00866e8c
36642006
09f260c3
0b84301c
0000311c
001c6c0c
3664211b
04c3988c
0100101c
08cb9cbc
4000201c
6126500e
a027702e
575c0894
61e64886
4006708e
00f350ae
575ca6f2
b08e4886
70ae61e6
6aac28c3
0483335c
7b8e78ce
1114301c
0000311c
6d2c6c0c
366406c3
0f568076
00000804
3f36f016
60c3fb96
92c3b1c3
cf5ca3c3
0f5c0203
00f70223
b830b80c
3bc3242b
301c4c4c
311c1114
6c0c0000
6c0c6c0c
03e3335c
4a946107
602774a9
000994dc
19e98500
0d940027
31e95a69
27d4301c
0015311c
259d333c
a4dc13e4
01330008
64dc0007
51e90008
23e47a69
000814dc
813791e9
1251365c
7a5434e4
0a940027
34c39a69
303c7fe5
765c300d
378309c4
00070173
1a696d94
5fe520c3
32236026
09a4165c
60073183
2f5c6394
265c0081
301c1255
311c1114
6c0c0000
04c4335c
15c306c3
366459e9
61a74013
79ec5194
0100093c
0260133c
eabc40c6
000708cb
74a94794
03546027
42946067
1110301c
0000311c
6e8c6c0c
20060086
70c33664
1114401c
0000411c
10940007
6c0c700c
21266c0c
03e6135c
a037700c
02868e4c
27c322a6
466437c3
40063a13
0456255c
59ec700c
06c36e6c
0260123c
366427c3
355c6026
e1c64ca6
03e6755c
6c0c700c
07e6735c
165c700c
013c1243
2fac3e87
301c4106
311c0b30
5abc0000
74a90874
50946027
4a41355c
4c946067
03e3355c
34dc6207
093c001a
153c0100
40c66ba0
08cbeabc
94dc0007
055c0019
30c349e1
0002341c
12546007
101c0186
111c0b30
b4bc0000
155c0873
21c349e1
00fd241c
3f5c40b7
355c0041
455c49e5
8ad24883
1114301c
0000311c
6e8c6c0c
200605c3
755c3664
e0074543
401c1254
411c1114
700c0000
06c36eac
701c2006
578008a8
700c3664
06c36ecc
36642006
055c0006
8a3c4a45
3c3c0240
73c3fdc0
06c37364
28c32546
d4bc37c3
40c30a88
602774a9
60670354
355c4294
620703e3
093c3e94
153c0100
40c66ba0
08cbeabc
35940007
33548007
31c33049
0002341c
0443255c
17946007
11544007
03f3255c
341c32c3
355cfffd
301c03f6
311c1114
6c0c0000
05c36eec
366416c3
355c6006
02730446
355c4ff2
617203f3
03f6355c
1114301c
0000311c
6eec6c0c
16c305c3
00263664
0446055c
00536046
54a96006
03544047
2a944007
0443255c
141c12c3
2077fffe
22942007
20548007
11a26045
341c30c3
60070001
1f5c1954
155c0021
4ff24ccd
03f3355c
355c6172
301c03f6
311c1114
6c0c0000
0dc36eec
366416c3
0443355c
355c6072
265c0446
40070989
06c31954
28c320e6
d4bc37c3
10c30a88
d2dc0007
6026000c
0ba5365c
1750063c
24c38429
b0bc4045
e00608cb
098d765c
355c17d3
620703e3
093c4694
153c0100
40c66ba0
08cbeabc
3d940007
602774a9
60670354
3bc33894
0683335c
455c7a6e
80073d19
701c1454
711c1114
7c0c0000
06c38f0c
60d718c3
5e8523c3
46646006
05d20364
6f2c7c0c
366406c3
455c8006
301c4526
311c1120
ec090000
1354e007
0c0d0006
1114301c
0000311c
055c6c0c
0a123653
41262fcc
0b30301c
0000311c
08745abc
03e3355c
47946207
0100093c
6ba0153c
eabc40c6
000708cb
79e93e94
3b946027
602774a9
60670354
44863694
323c0653
1ac30010
60090580
24a72522
155c2694
60094a16
351c6812
355c0025
323c4a16
33640020
5da27ac3
4a26255c
04293d80
412c303c
4a26355c
255c4449
60264a35
4a45355c
1114301c
0000311c
6f4c6c0c
202606c3
06333664
69806045
236423c3
ce142ce4
03e3355c
1d946207
0100093c
6ba0153c
eabc40c6
000708cb
79e91494
11946027
002714a9
00670354
301c0c94
311c1114
6c0c0000
06c36f6c
2cc31ac3
0bf23664
105c201c
0000211c
34c3880b
680e6025
00530006
05960026
0f56fc76
00000804
0f36f016
61c3fe96
a3c392c3
a00ca364
2f5c4006
6a06002d
00353f5c
1f5c3e46
8006003d
0050bf3c
fa000953
0009875c
331c7a22
3e9400dd
0020343c
1bc31980
2abc4066
01640892
34940007
60477ca9
74a93194
03546027
24946067
3d19255c
355c4ad2
5a003481
21c32909
000f241c
205432e4
4d097a00
341c32c3
6037000f
00013f5c
3485355c
00a0343c
6800053c
42063980
08cbb0bc
155c2026
00263d1d
3a3c0233
540c05c7
20266d00
0175135c
383c0133
71800020
436443c3
b67449e4
02960006
0f56f076
00000804
0336f016
80c3fc96
12c361c3
73c31264
5f5c7164
0f5c0161
00770181
880c28c3
402749e9
153c2494
2037fcc0
00013f5c
19b46b07
30c3192b
0100341c
13946007
39222213
6c297900
b2dc24a7
42870010
24f20594
52dc6007
60450010
23c36980
00532364
27e44286
03b3ed74
32a331c3
60072286
02f31654
788058a2
40670c29
6c490594
085435e4
22871d93
44f20594
72dc0007
303c000e
65800020
136413c3
eb7417e4
0440783c
0ebc07c3
01640892
1aa900f7
301c00b7
311c0ba0
2c0b0000
341c31c3
60070040
301c1154
311c1114
6c0c0000
0604535c
06c3a9d2
00212f5c
400612c3
0160363c
08c35664
0359105c
341c31c3
60070001
545c2c54
a10703e3
305c2894
600707d3
00972494
00d710c3
1f9410e4
0160063c
3f5c17c3
23c30041
08922abc
00070164
301c1494
311c1114
6c0c0000
6c0c6c0c
035c0126
05c303e6
0b30101c
0000111c
0873b4bc
11930046
03e3345c
0e946207
602770a9
345c0bb4
68d24543
08e8101c
0ebc1080
01640892
40d700f7
600732c3
70a976f4
07946067
0160063c
3f5c17c3
09b30061
03e3345c
11b461e7
10c30097
10e400d7
063c6294
17c30160
00413f5c
2abc23c3
01640892
57940007
03e3345c
1e946207
602770a9
145c1b94
20074543
245c1754
400745b1
60971394
60d793c3
439493e4
0160063c
08e8201c
3f5c3100
23c30041
08922abc
00070164
345c3694
620703e3
10a91a94
17940007
4543145c
13542007
32c34097
32e440d7
063c2694
301c0160
318008e8
00413f5c
2abc23c3
01640892
19940007
03e3345c
17b461e7
10c30097
10e400d7
063c1294
17c30160
00413f5c
2abc23c3
01640892
202608f2
105c08c3
00730835
00531fe6
04960026
0f56c076
00000804
ff963016
301c40c3
311c1114
0c0c0000
508c202c
67d26849
341c680c
331cf000
0c945000
6c0c600c
50c30929
503c0c89
a03732ac
00013f5c
680c692d
f000341c
29946007
78bc0106
201c08cc
211c0bb4
325c0000
602507a4
07a7325c
07e4325c
425c64f2
005307c7
301c8c0f
311c0bb4
435c0000
a00607e7
0106b00f
08cc82bc
15c300a6
0fe4301c
0000311c
d4bc4d0c
02d308c8
6025640c
644c640f
842f63f2
8c0f0053
0006844f
301c100f
311c1114
6c0c0000
135c6c4c
a2bc1341
01960872
08040c56
51c37016
600c5364
48e4435c
1101245c
354332c3
0014633c
1e94c007
1114301c
0000311c
6dec6c0c
36640026
0247153c
fc7f301c
000a311c
02e423c3
70800ab4
3500201c
000c211c
235c4820
00930b47
635c7080
0e560b47
00000804
30c3ff96
60873264
60a70514
60e70635
60060735
01336037
3444315c
315c0073
233c3464
4037090b
00013f5c
019603c3
00000804
fe967016
533c608c
8c890100
61891600
1d946107
600761a9
615c1a94
c0073d19
301c1254
311c1114
6c0c0000
053201e9
335c0037
2f5c05a4
02c30001
30c33664
65f23264
6de97600
00536532
60776006
00216f5c
029606c3
08040e56
0736f016
70c3f596
427791c3
2109c00c
42d223d2
29c3c02c
a55ca88c
22570021
05c7313c
6d00580c
0223135c
746c2fd2
211c4006
3283000f
111c2006
21c3000b
045432e4
8000301c
301c74ce
311c1114
6c0c0000
09c36d0c
366416c3
326430c3
23c362b7
42375fe5
01013f5c
1c356027
43d24297
04944067
0001801c
229702f3
5f8521c3
3f5c41f7
801c00e1
60270002
42970d35
7f4532c3
3f5c61b7
801c00c1
60270003
801c0335
78a90000
03546047
14946007
1114301c
0000311c
1f5c6c0c
1f5c0141
8f5c0005
435c0027
07c30524
425719c3
466436c3
275c1b73
47d203a1
74cd6026
6c0c7c0c
348e2feb
40067dac
0008211c
60073283
365c3054
620703e3
265c2c94
40073d19
365c2854
60073d09
265c2454
682b48e4
1fb46027
31c32257
61126145
4c2b6980
429732c3
233c3243
40070014
301c1294
311c1114
6c0c0000
1f5c2f89
22570005
00261f5c
07c38d4c
13c36297
46646046
383c746c
2297241b
251b313c
2f5c746f
55ed0121
3d19365c
74cb64d2
74ce6c72
01c0353c
4c801ac3
49a3365c
37546007
331c6809
33940088
331c6829
2f94008e
29c36086
01d5325c
4086740c
231b323c
2006740f
5469344d
500632c3
617732a3
00a13f5c
301c746d
311c1114
6c0c0000
0544435c
15c307c3
602626c3
35294664
241c21c3
413700c0
00813f5c
35c3752d
033e133c
241c21c3
08b3fdff
03e3365c
42946207
331c6809
3e940088
331c6829
3a94008e
1114301c
0000311c
435c6c0c
07c30544
26c315c3
46646026
13c37529
00c0141c
2f5c20f7
552d0061
39c32086
01d5135c
4086740c
231b323c
4006740f
7469544d
700613c3
20b713a3
00411f5c
35c3346d
033e133c
241c21c3
4c0efdff
4d89265c
35c349f2
063e133c
101c21c3
21a38000
301c4c0e
311c1114
6c0c0000
09c36d2c
00063664
e0760b96
08040f56
3f36f016
0277ee96
52c391c3
435c600c
21c348e4
0980642b
61004089
82c34e09
0001841c
600738c3
80304694
40063cc3
0100211c
60073283
61c93e54
241c23c3
4107000f
353c38b4
043c0020
30c3359d
341c3263
60070001
353c2e54
6d00180c
743c6285
e067359d
373c26b4
71800247
14c0233c
0003b25c
4377482b
0a83635c
0a53a35c
0b23d35c
630bcc3c
84dccbe4
6026000a
700d133c
2f5c2437
42b70201
023702e3
01011f5c
573c22f7
ca3c0097
07d3fff0
1114301c
0000311c
6dcc6c0c
366409c3
245c3c93
04171101
328330c3
6de46bd2
62d70994
028303c3
1f5c01f7
145c00e1
201c1105
211c1114
680c0000
09c36dcc
383c3664
83c30010
77008364
20066aa5
3b9d143c
00103b3c
fff4b33c
32c34357
133c6025
2377fff4
0010363c
63c33c83
77006364
943c6aa5
29c33a1d
ca944007
0001831c
0019d9dc
1101045c
374330c3
0001341c
44dc6007
56c30019
0097c73c
fff09a3c
1cc30813
6aa56680
3a1d343c
30546007
1101245c
30c30417
d5c33283
28946007
101c4bd2
111c1114
640c0000
02576e0c
366417c3
201c0253
211c1114
680c0000
0800001c
2faf011c
41462fec
0b30301c
0000311c
08745abc
03c36297
1101345c
01b703a3
00c10f5c
1105045c
353cd5c3
39830010
536453c3
0010383c
836483c3
c0948ae4
2cc32973
323c2ba4
3ae4fff4
79005315
fff02a3c
53c33283
373c5364
6e800097
343c6aa5
60073a1d
301c1154
311c1114
6c0c0000
6c6c6c4c
05a4235c
0bb4301c
0000311c
26640c0c
245c2693
323c1101
341c708d
60070001
301c2694
311c1114
47d20000
6e0c6c0c
17c30257
01d33664
001c6c0c
011c0800
2fec2faf
301c4146
311c0b30
5abc0000
60260874
700d233c
345c4177
23a31101
0f5c4177
045c00a1
d5c31105
0097373c
6aa56e80
3b9d943c
323c1e73
331cfff4
c6dc0800
3cc3000d
321c3aa4
233c1001
4337fff4
133c6026
2477700d
02212f5c
02e343b7
1f5c0137
23f70081
0097373c
1a3c6077
2037fff0
40570693
533c6b00
043c0550
0bd25a1d
1114101c
0000111c
6dcc640c
40063664
5b9d243c
1101245c
30c30457
6bd23283
09946de4
03c363d7
00f70283
00611f5c
1105145c
0010383c
836483c3
00103b3c
fff4b33c
03948ae4
0173c006
0010363c
30830017
636463c3
21c32317
ca94b2e4
fff03a3c
4f003364
a164a3c3
528353c3
0097273c
6aa56a80
3b9d943c
01a7cf5c
31c32317
4094b3e4
6aa56b00
3a1d043c
01a7cf5c
1114901c
0000911c
065382c3
640c19c3
36646dcc
1101245c
30c30457
6bd23283
09946de4
03c363d7
00b70283
00411f5c
1105145c
6b0028c3
00066aa5
3b9d043c
0010363c
23832ac3
636462c3
30c30317
233c6025
4337fff4
30c30357
233c6025
4377fff4
630008c3
043c6aa5
00073a1d
245cce94
323c1101
341c708d
60070001
373c3f94
6e800097
343c6aa5
60073a1d
301c3754
311c1114
47d20000
6e0c6c0c
17c30257
01d33664
001c6c0c
011c0800
2fec2faf
301c4146
311c0b30
5abc0000
23970874
145c21c3
21a31101
2f5c43b7
245c01c1
bf5c1105
d5c30184
301c0273
311c1114
6c0c0000
6c6c6c4c
05a4235c
0bb4301c
0000311c
26640c0c
bf5c0073
373c0184
71800247
14c0233c
0006b25c
082e0357
0a86635c
0b26d35c
fc761296
08040f56
50c33016
301c5364
311c1114
6c0c0000
52098c8c
354332c3
0001341c
00c66ad2
089580bc
5a1d343c
031c0180
02b407cf
0c560006
00000804
0136f016
81c370c3
026402c3
5d09dc0c
02d243d2
380cdc2c
8c0938c3
241c24c3
40070001
78a92094
06546027
05c0413c
606752c3
00061394
043c02d3
18c30010
eabc40c6
08f208cb
033c7009
9d090010
03c38ad2
8b850113
365ca025
53e403a3
1fe6ed14
0f568076
00000804
6e676962
655f6d75
6d747078
685f646f
00000077
70797263
6d5f6f74
655f646f
685f7078
00000077
636c6163
5f68645f
0079656b
4d5f4e4e
0000646f
00240000
002c0028
00340030
003c0038
00640040
006c0068
00740070
007c0078
00840080
008c0088
00990095
00a1009d
000000a5
103c1016
203cb80b
403c45cb
0006f88c
18f44fc7
ffff301c
7fff311c
231c1180
10d4009d
177201c3
0095231c
323c05f4
0323f6a0
301c00b3
6d200096
82d20343
085600c4
00000804
20c37016
200630c3
ffff111c
333c3183
7fe50b0d
633c7f32
6206200c
23636f20
341c32c3
7fe5ff00
533c7f32
6106180c
23636ea0
0f04323c
7f327fe5
100c433c
6e206086
310d123c
00c4313c
7f327fe5
080c233c
61200046
77001363
8d006e00
0026313c
084b333c
40a033c4
11803283
08040e56
20c31016
000710c3
101c3754
131c009e
0ef40099
301c0006
6ca000b9
300d323c
002662d2
f670313c
308d323c
301c03a3
4ca00099
400730c3
303c03f4
23c3200d
341c5a92
6087000f
40850254
800632c3
0400411c
69d23483
313c5a92
333c0fe6
33c40b0d
23837f52
101c4332
44d200ff
101c5672
600600ff
b81b323c
45db313c
03c37f92
08040856
03f27016
0b9301c3
200751c3
103c5954
653c45cb
363c45cb
13e40190
313c51d4
63e40190
05c303f4
30c30973
ffff201c
007f211c
77723283
300c433c
328335c3
233c7772
0007300c
44c40215
0215a007
16e422c4
672004f4
00932363
436378a0
4a0016c3
06154007
800622c4
8000411c
000600f3
44f240c3
41120473
32c33fe5
011c0006
3083e000
32c379d2
011c0006
30834000
415263d2
323c2025
63e5098b
32c34d00
011c0006
30834000
415263d2
323c2025
013c310c
7792ba2c
0e5603a3
00000804
21c330c3
06f22ed2
111c2006
68808000
60060113
8000311c
a6bc2580
30c30a94
080403c3
000730c3
20070815
40060615
8000211c
25006100
31e41fe6
00060574
02f431e4
08040026
0336f016
03d260c3
23f251c3
09b30006
45cb203c
45cb313c
938492c3
f820793c
201c30c3
211cffff
3283007f
377213c3
328335c3
177203c3
410c413c
410c203c
428d823c
0ff4313c
228d333c
410c233c
0ff4303c
428d333c
69806852
233c3884
32c3108c
111c2006
31832000
323c66d2
233c0200
00f3308c
0100323c
288c233c
f810793c
200632c3
0100111c
63d23183
e0254132
60066503
8000311c
073c6383
32c3bb2c
03a37792
0f56c076
00000804
60c3f016
40066103
8000211c
2af26283
211c4006
c0074f80
40063794
4f00211c
20c30673
30540007
45cb303c
07e0233c
45cb313c
30c3a9a0
ffff701c
007f711c
03c33783
17831772
977241c3
031504e4
bfe50112
20064006
0100111c
04e432c3
21a30374
01120220
60252152
f8946327
0010323c
090c133c
0010353c
bb2c233c
779231c3
02c323a3
08040f56
05d230c3
211c4006
61008000
080403c3
20c3fe96
605703f2
600665d2
8000311c
02c34180
08040296
30c3fe96
203c0fd2
30c3a0cb
111c2006
31838000
303c23a3
321c45cb
333c0380
03c3a12c
08040296
05f2fe96
23c36057
1d546007
5d0b303c
c800133c
201c30c3
211cffff
3283000f
547223c3
76326057
51ac323c
60256632
77926152
b9ac313c
211c4006
02838000
20a323c3
029602c3
00000804
00b7fc96
00072037
20070a15
40060815
8000211c
60b76100
60376500
60174097
0d7423e4
23e40026
40d70bd4
23e46057
00060614
043523e4
00530026
04961fe6
00000804
fe963016
04f210c3
60076057
413c2954
543c5d0b
0057be30
0bf4a007
011c0006
20078000
001c1e74
011cffff
03337fff
201c31c3
211cffff
3283000f
547223c3
b08c303c
51ac023c
c020343c
08b463c7
35c407d2
20070363
00c40415
00060053
0c560296
00000804
fe963016
003740c3
605704f2
2d546007
5d0b343c
bc20233c
20570017
0df44007
20060006
8000111c
217440e4
101c1fe6
111cffff
03737fff
fc01321c
15b467c7
ffff301c
000f311c
34721383
e0bc22c4
20c30a7c
800731c3
02c40a15
02f22026
33c410c3
00732ca0
10c30006
0c560296
00000804
fe963016
04f210c3
60076057
413c1b54
543c5d0b
4057be20
a0071fe6
301c14d4
311cffff
1383000f
747231c3
033c5532
343c592c
63c7c010
04d205b4
034335c4
00060053
0c560296
00000804
fe967016
30c3a057
600735a3
203c1354
423c5d0b
7fe6bc20
800713c3
323c0dd4
67c7c010
15c307b4
a4bc24c4
30c30a7c
60060073
03c313c3
0e560296
00000804
0336f016
00b7fc96
31c38057
600734a3
000982dc
30c340d7
6ed232a3
5d0b903c
5d0b813c
0360383c
b6dc93e4
393c0008
83e40360
20b703f4
301c1093
311cffff
2383000f
303c5472
723cb88c
503c49ac
201c480c
211cffff
4283000f
547224c3
b88c313c
49ac623c
480c413c
08150007
402605c4
20c302f2
50c337c4
2007ed20
04c40815
02f24026
36c420c3
cd2040c3
0af498e4
16c304c3
28a429c3
0a7ce0bc
61c340c3
05c30133
28c317c3
e0bc29a4
50c30a7c
528071c3
24e42026
20060214
65807b80
13c302c3
05746007
31a332c3
06d36ef2
202602c4
10c302f2
2ca033c4
303c00d3
0112f88c
09ac113c
a00631c3
e000511c
76d23583
400631c3
c000211c
65d23283
013c0132
2152f82c
0a4b303c
00ff321c
40260c00
021403e4
28804006
a00631c3
c000511c
66d23583
088c303c
f9ac013c
303c2152
313c488c
60b7b9ac
04960097
0f56c076
00000804
fc961016
31c320c3
34a38057
40066fd2
8000211c
20372500
00b730c3
34a380d7
64d221c3
0a96eebc
02c320c3
08560496
00000804
0f36f016
80c3fc96
38c300d7
66d230a3
405791c3
32a331c3
a00664f2
1013a0b7
ffff101c
000f111c
30c30183
21837472
583c5472
533ca88c
733c5aac
493ca90c
423ca88c
623c5a2c
04c3a90c
25c316c3
5abc37c3
a0c30a7e
08c3b1c3
ffff101c
001f111c
20060183
36c324c3
0a7e5abc
a88c403c
5a2c413c
a90c613c
201c09c3
211cffff
0283001f
25c32006
5abc37c3
303c0a7e
313ca88c
355259ac
4026b180
021454e4
78804006
4ac34980
20261600
021405e4
4bc32006
65806a00
033c0232
233cf02c
32c3108c
511ca006
35832000
403c6fd2
20261000
021440e4
65002006
488c043c
b82c033c
488c133c
403c01d3
20260800
021440e4
650013c3
408c043c
c02c033c
408c133c
400631c3
0020211c
65d23283
088c303c
f9ac013c
009700b7
f0760496
08040f56
0f36f016
b1c3fc96
20c360d7
205723a3
3bc347f2
67f231a3
20b73fe6
2bc30b33
43f221a3
0a9340b7
ffff201c
000f211c
23c33283
00b75472
301c40f7
311cffff
1383000f
91c33472
05d412e4
0b9492e4
0935b0e4
f88c303c
09ac223c
080c303c
40f760b7
20d74097
c0060006
0020611c
a0c370c3
91e480c3
91e411d4
b2e40394
70a30db4
3bc3a6a3
8026a9a0
02b452e4
29c38006
25c36520
323c2e20
4112f88c
09ac113c
088c303c
f9ac063c
821cc152
831c0001
e0940036
0010373c
37e44026
40060214
61322a84
f9ac323c
009760b7
f0760496
08040f56
0a9618bc
f90c303c
033c6c20
0804f88c
0a951abc
f90c303c
033c6c20
0804f88c
0a9618bc
08041f52
0a951abc
08041f52
0a9618bc
08041f52
0a951abc
08041f52
0a9618bc
f90c303c
033c6c20
0804f88c
0a951abc
f90c303c
033c6c20
0804f88c
fe961016
21c30077
30c32006
089432e4
3fc34097
04c38c2c
029420e4
01c32026
08560296
00000804
21c3fe96
30c32006
029432e4
01c32026
08040296
fe961016
21c30077
30c32006
079432e4
3fc34097
04c38c2c
025420e4
01c32026
08560296
00000804
21c3fe96
30c32006
025432e4
01c32026
08040296
001c30c3
64d2ff53
0967135c
08040006
61e6fe96
21c321a2
40374025
00011f5c
2f5c2077
41a10021
7fe524f2
f3947fe7
08040296
61e6fe96
21c321a2
40374025
00011f5c
2f5c2077
41a10021
7fe524f2
f3946167
08040296
3f36f016
a0c3fb96
e00c2137
2ac3c02c
044e123c
082c82c3
a077a006
a0b7a0f7
411795c3
398432c3
40374c0c
c01cac30
d31c0000
0e150000
32c340d7
60f73703
32c34097
60b73603
40575103
300332c3
313c6077
273c0014
60070014
80061a54
8000411c
800642f2
088c313c
088c203c
f9ac103c
02a304c3
088c373c
088c263c
f9ac763c
600662c3
e100311c
02d36303
8006b3c3
8000411c
43c342f2
088c313c
f9ac303c
088c203c
13a31bc3
02a304c3
088c373c
f9ac763c
c21cc132
c31c0001
09540040
7f326017
41124017
dd3c4037
f61309ac
0008921c
0010931c
60d7a394
680f2ac3
682f6097
a80f28c3
682f6057
fc760596
08040f56
fe961016
01d36006
42c341e9
80378025
00012f5c
4f5c4077
81ed0021
44f21fe5
31e46025
0296f214
08040856
60c37016
43c352c3
b0bc25d2
565c08cb
87d208a7
0f40063c
420614c3
08cbb0bc
0e560006
00000804
ff961016
803780d7
0a99d8bc
08560196
00000804
ff961016
06544207
04544307
09944407
44070073
80d706b4
d8bc8037
00730a99
ff53001c
08560196
00000804
fb96f016
71c360c3
420752c3
43070554
44070354
4f3c1094
04c30040
42062006
0891b0bc
60376006
17c306c3
34c325c3
0a99f6bc
0f560596
00000804
30c3ff96
001c2037
6007ff53
033c1154
60170f40
420666d2
08cbb0bc
01130006
00013f5c
420613c3
0891b0bc
01960017
00000804
3f36f016
40c3f296
92c361c3
df5cc3c3
bf3c0324
0bc30280
4c84101c
0016111c
e6bc4206
5f3c08cb
05c30180
1180143c
b0bc4206
05c308cb
420615c3
0b0672bc
200719c3
c0076254
893c6054
a93c208c
46c300f4
00078f5c
00807f3c
07c30493
420614c3
08cbb0bc
17c307c3
72bc4206
60970b06
229740d7
22d73103
62b72103
611742f7
23174157
23573103
63372103
0bc34377
46bc15c3
82050a99
32c34017
60377fe5
20072017
383cdb94
b980200c
40072ac3
4f3c2a54
04c30080
00013f5c
420613c3
0891b0bc
15c304c3
b0bc2ac3
04c308cb
420614c3
0b0672bc
40d76097
31032297
210322d7
42f762b7
41576117
31032317
21032357
43776337
02800f3c
01801f3c
0a9946bc
40072dc3
3cc36654
63546007
208c6d3c
00f47d3c
c0774cc3
00805f3c
0280af3c
01808f3c
05c30493
420614c3
08cbb0bc
15c305c3
72bc4206
60970b06
229740d7
22d73103
62b72103
611742f7
23174157
23573103
63372103
0ac34377
46bc18c3
82050a99
32c34057
60777fe5
20072057
363cdb94
2cc3200c
e007a980
4f3c2a54
04c30080
00213f5c
420613c3
0891b0bc
15c304c3
b0bc27c3
04c308cb
420614c3
0b0672bc
40d76097
31032297
210322d7
42f762b7
41576117
31032317
21032357
43776337
02800f3c
01801f3c
0a9946bc
e88c293c
393c6297
22d7199c
62b72103
2d3c42f7
6317e88c
199c3d3c
21032357
43776337
02804f3c
1f3c04c3
46bc0180
04c30a99
420614c3
0b0672bc
14c30697
b0bc46d7
0e9608cb
0f56fc76
00000804
0336f016
50c3fd96
72c391c3
305c83c3
400608a4
620740b7
361c0b54
333c0018
7fe50b0d
f88c233c
6d206046
653c60b7
383c1040
06c3ff00
42063d80
08cbb0bc
f5248e24
78bc0126
05c308cc
00413f5c
54bc13c3
053c087c
2f5c0f40
12c30041
087c88bc
00413f5c
00053f5c
00279f5c
18c307c3
60064026
087cbcbc
82bc0126
343c08cc
62d24004
053cf324
16c30f40
b0bc4206
000608cb
c0760396
08040f56
0336f016
70c3fd96
82c391c3
305c63c3
400608a4
620740b7
361c0b54
333c0018
7fe50b0d
f88c233c
6d206046
301c60b7
311c10f8
6c0c0000
06c38c0c
44c62006
4c94301c
0016311c
50c34664
26c318c3
08cbb0bc
f5248e24
78bc0126
07c308cc
00413f5c
54bc13c3
073c087c
2f5c0f40
12c30041
087c88bc
00413f5c
00053f5c
05c3a077
400616c3
bcbc32c3
0126087c
08cc82bc
4004343c
f32462d2
ff00363c
0f40073c
42063580
08cbb0bc
15c309c3
b0bc26c3
301c08cb
311c10f8
6c0c0000
05c38c4c
44c62006
4c94301c
0016311c
00064664
c0760396
08040f56
fd96f016
61c350c3
305c72c3
400608a4
620740b7
361c0b54
333c0018
7fe50b0d
f88c233c
6d206046
053c60b7
16c31040
b0bc4206
8e2408cb
0126f524
08cc78bc
3f5c05c3
13c30041
087c54bc
00412f5c
00052f5c
06c3e077
40262206
bcbc32c3
0126087c
08cc82bc
4004343c
f32462d2
0f560396
00000804
12c331c3
16bc23c3
08040a9c
0136f016
60c3fd96
82c371c3
08a4305c
40b74006
0b546207
0018361c
0b0d333c
233c7fe5
6046f88c
60b76d20
10f8301c
0000311c
8c0c6c0c
20060206
301c44c6
311c4ca8
46640016
000750c3
17c33554
b0bc4206
8e2408cb
0126f524
08cc78bc
3f5c06c3
13c30041
087c54bc
00412f5c
00052f5c
05c3a077
40062206
bcbc6026
0126087c
08cc82bc
4004343c
f32462d2
15c308c3
b0bc4206
301c08cb
311c10f8
6c0c0000
05c38c4c
44c62006
4ca8301c
0016311c
03964664
0f568076
00000804
0336f016
81c390c3
63c372c3
42c351c3
06c301b3
420615c3
0b0696bc
9e05a205
16c309c3
58bc26c3
81e70a9c
37c3f3b4
32835e06
08c35da0
49d22180
96bc06c3
09c30b06
26c316c3
0a9c58bc
0f56c076
00000804
0136f016
80c3f896
52c371c3
12c363c3
ff00141c
009f233c
feff001c
0000011c
54e440c3
413c11b4
4203408c
1f5c81f7
380d00e1
4c0945c3
81b74203
00c14f5c
00468c0d
42e30733
0f5c8177
180d00a1
42c34c09
42035fc6
4f5c8137
8c0d0081
253c36c3
40f7c08c
011e433c
40f72403
00610f5c
36c30c0d
440b453c
033c80b7
4003019e
2f5c80b7
4c0d0041
013c36c3
0077408c
021e133c
00770103
00212f5c
36c34c0d
433c05c3
0403029e
0f5c0037
0c0d0001
620600c6
18008c20
081454e4
24c317c3
0b0696bc
fe00b620
17c300d3
96bc25c3
a0060b06
16c308c3
58bc26c3
a7d20a9c
17c308c3
36c325c3
0a9cb8bc
80760896
08040f56
3f36f016
80c3f196
c2c32137
269793c3
000786d7
001002dc
40074117
000fc2dc
60073cc3
000f82dc
52dc2007
a717000f
12dca007
80c7000f
000ee9dc
b5dc81a7
0f3c000e
24c301d0
08cbb0bc
6e2061e6
4f5c60f7
81b70061
80b79fe5
00411f5c
2f5c2177
2f5c00a1
6f3c00e5
d6c302b0
7a208197
200600f3
d21c5dc3
153cffff
d3e4ffdf
6026f994
015d3f5c
800659c3
02c0af3c
08c302f3
01c01f3c
58bc2ac3
0ac30a9c
420617c3
0b0696bc
1ac30bc3
b0bc4206
0f3c08cb
219701c0
0a99c2bc
2117be05
b484b1c3
ea002cc3
a1e78205
39c3e3b4
34839e06
f5a059c3
a384a1c3
29c3a980
13544007
02c04f3c
1f3c08c3
24c301c0
0a9c58bc
15c304c3
96bc27c3
0ac30b06
27c314c3
08cbb0bc
009336c3
433c8006
3de4ffdf
08c3fc94
01c01f3c
02c02f3c
0a9c58bc
47d72806
12c342f2
03a13f5c
ffe0233c
f88c323c
61526d00
81576312
65807180
5f5c6077
5f5c0021
06c300e5
101c4006
24d200ff
02354067
323c2006
393c18dc
51c3308d
a0375383
00013f5c
ffdf303c
81974025
25e454c3
4f3ced14
08c302c0
01c01f3c
58bc24c3
27d70a9c
08c327d2
47d72797
e2bc34c3
29c30a9c
08c347d2
3f3c2117
b8bc02c0
3f5c0a9c
3f5c00a1
009300e5
463c8006
6de4ffdf
4f3cfc94
08c301c0
24c314c3
0a9c58bc
02c05f3c
14c305c3
96bc4757
05c30b06
47572717
0b06c0bc
08d240c3
20060117
b0bc29c3
401c0891
0f3cff4b
220602c0
0b06b8bc
01c00f3c
b8bc2206
00730b06
ff53401c
0f9604c3
0f56fc76
00000804
3f36f016
80c3f396
c2c3d1c3
2617a3c3
e6978657
0007c757
000da2dc
40072dc3
000d62dc
60073cc3
000d22dc
f2dc2007
e007000c
000cc2dc
99dc80c7
81a7000c
000c65dc
01500f3c
b0bc24c3
61e608cb
60f76e20
00612f5c
b264b2c3
c2f22806
5b3c16c3
a0b7fff0
00412f5c
3f5c4137
233c0361
323cffe0
6d00f88c
63126152
7580a117
60776580
00212f5c
00a52f5c
02304f3c
400604c3
00ff101c
24d20253
02354067
323c2006
3a3c18dc
91c3308d
9f5c9383
3f5c0007
303c0001
4025ffdf
ee142be4
02405f3c
1f3c08c3
25c30140
0a9c58bc
08c3c7d2
26c32717
e2bc35c3
2ac30a9c
08c347d2
3f3c1cc3
b8bc0240
07c30a9c
02401f3c
b0bc46d7
5f3c08cb
3f5c0340
353c0081
3f3cf05e
3ba40230
40060093
ffdf243c
fc9443e4
02404f3c
15c308c3
58bc24c3
07c30a9c
46d714c3
0b0696bc
2f5c4026
7ac3011d
02f3c006
1f3c08c3
24c30140
0a9c58bc
15c304c3
96bc4206
09c30b06
420614c3
08cbb0bc
01400f3c
c2bc1bc3
fe050a99
96849dc3
ab002cc3
e1e7c205
3ac3e4b4
3583be06
a9a02ac3
c9802cc3
e9802dc3
1354a007
02404f3c
1f3c08c3
24c30140
0a9c58bc
16c304c3
96bc25c3
07c30b06
25c314c3
08cbb0bc
02400f3c
b8bc2206
0f3c0b06
22060140
0b06b8bc
00730006
ff53001c
fc760d96
08040f56
3f36f016
90c3e896
b2c320f7
c8d7c3c3
4f3ca917
04c30400
42062006
0891b0bc
0a94a187
16c304c3
b0bc25c3
602608cb
027d3f5c
a0370173
42068077
09c340b7
21c32006
44bc36c3
6f3c0a9a
06c30500
04001f3c
b0bc4206
cf5c08cb
5f3c0007
a0770200
60b76206
29d709c3
3bc34a17
0a9a44bc
01004f3c
16c309c3
58bc24c3
05c30a9c
420614c3
0b0696bc
15c30957
c0bc4997
30c30b06
ff4c001c
46946007
208cac3c
43c37ac3
5f3cd6c3
02930300
34bc0dc3
09c30a99
25c31dc3
0a9c58bc
16c305c3
96bc4206
08c30b06
420615c3
08cbb0bc
40d7ffe5
848482c3
ce003bc3
e0078205
3a3ce694
a2c3200c
8bc3a384
6c3c8384
07c300f4
1854c007
05005f3c
34bc05c3
4f3c0a99
09c30300
24c315c3
0a9c58bc
18c304c3
96bc26c3
0ac30b06
26c314c3
08cbb0bc
189607c3
0f56fc76
00000804
3f36f016
90c3f096
40f7d1c3
c6d7b3c3
a33ca717
4f3c00f4
04c30200
42062006
0891b0bc
0a94a187
16c304c3
b0bc25c3
602608cb
017d3f5c
a0370173
42068077
09c340b7
21c32006
44bc36c3
cb3c0a9a
4f3c208c
04c30300
02001f3c
b0bc4206
6cc308cb
4f3ca006
02d30100
03000f3c
0a9934bc
1f3c09c3
24c30300
0a9c58bc
17c304c3
96bc4206
08c30b06
420614c3
08cbb0bc
8dc3dfe5
40d78584
a205ea80
e594c007
200c3c3c
e9802dc3
c98040d7
60073ac3
5f3c1754
05c30300
0a9934bc
01004f3c
15c309c3
58bc24c3
04c30a9c
2ac316c3
0b0696bc
14c307c3
b0bc2ac3
bf5c08cb
47570007
67974077
09c360b7
481727d7
44bc3dc3
4f3c0a9a
09c30100
02001f3c
58bc24c3
07570a9c
479714c3
0b0696bc
10960006
0f56fc76
00000804
2037fa96
42174077
425740b7
613740f7
617761d7
21c32006
f6bc31c3
06960a9f
00000804
0136f016
70c3fb96
52c381c3
07544207
05544307
ff53401c
18944407
00406f3c
200606c3
b0bc4206
60060891
07c36037
25c318c3
f6bc36c3
40c30a99
07c307f2
273c16c3
58bc1180
04c30a9c
80760596
08040f56
0aa098bc
00000804
3f36f016
40c3fe96
92c3a1c3
c03c53c3
0cc31040
0944145c
133c60a0
03130100
009f213c
921c69c3
363c0001
62c3009f
c0776303
00212f5c
a21c0ac3
203c0001
345c00df
7fe50944
0947345c
345cbfe5
63d20944
e594a007
743cd5c3
c0060f40
04c30253
28c317c3
0a9c58bc
22bc07c3
08c30a99
42061bc3
0b0696bc
6006be05
0947345c
b684b9c3
86848ac3
a1e7c205
3dc3e9b4
3683de06
a1a00dc3
838489c3
c9802ac3
2154a007
17c304c3
58bc2cc3
07c30a9c
0a9922bc
345c6206
40060947
21220cc3
08c331c3
01c32122
60373003
00011f5c
345c3921
7fe50944
0947345c
bfe54025
ed94a007
fc760296
08040f56
12c331c3
58bc23c3
08040a9c
0336f016
50c3fe96
92c371c3
400d4026
602d6006
80778006
7700c057
00212f5c
c0254c4d
631cc077
f7940100
01c32006
548041c3
c037c849
868484c3
dc2248c3
433c7300
76000ff4
011e633c
2f5cc84d
4c0d0001
09e40025
00060214
131c2025
e8940100
c0760296
08040f56
fd963016
69a2600c
840c6077
341c6e00
640f00ff
60b769a2
5f5c600c
a9a10041
1f5c640c
29a10021
43c36009
80378025
00015f5c
0097a00f
60802057
00ff341c
039609a2
08040c56
0f36f016
50c3fd96
82c391c3
400963c3
602940b7
703c6077
80060020
0080bf3c
0040af3c
28c30273
40374a22
1ac30bc3
7abc27c3
60170aa1
200323c3
2f5c4037
39c30001
80254e21
c007dfe5
3f5ced94
740d0041
00212f5c
0396542d
0f56f076
00000804
326430c3
fd00033c
00000804
0136f016
61c350c3
680c82c3
0010733c
d0bc05a2
303c0aa1
540c00a7
940f8d00
d0bc1ba2
70000aa1
373c740f
28c30010
8076680f
08040f56
ff96f016
61c350c3
43c372c3
4006040c
103c5c0f
14e40010
54001fb4
a037a809
00013f5c
05c33064
0e156007
07f4303c
00062580
063514e4
a80901f3
42ac003c
40257fe5
60807bf2
06b434e4
0007380f
1c0f05f4
001c0073
0196ff7c
08040f56
fe967016
52c341c3
40775fe6
2037240c
460740a2
213c1494
1f3c0010
213c0080
1fc3fc7e
00402f3c
0aa1f2bc
07740007
740f6057
d00fc017
007303c3
ff74001c
0e560296
00000804
fe967016
52c341c3
40775fe6
2037240c
462740a2
213c1494
1f3c0010
213c0080
1fc3fc7e
00402f3c
0aa1f2bc
07740007
740f6057
d00fc017
007303c3
ff74001c
0e560296
00000804
40c37016
440c52c3
001c6122
6047ff74
40250e94
001c7122
6027ff73
323c0894
91a20010
6025940f
140c640f
08040e56
61c3f016
440c42c3
700f6006
64092100
16946047
0010523c
20c302a2
08350087
700c01f3
333ce429
700f43ac
20255fe5
353c59f2
6c000010
100c780f
001c0073
0f56ff74
00000804
840cf016
331c6222
079400a0
0020343c
6abc640f
00930aa2
680f6006
0f5603c3
00000804
ff967016
62c351c3
41a2640c
640f6025
ff70401c
0e9440c7
36c32fc3
0aa1f2bc
ff74401c
06740007
4017740c
740f6d00
04c38006
0e560196
00000804
40c33016
ff7b001c
a0a6080f
8027ac0f
20271094
20670454
00d32194
280f2066
4c0f4186
a04601d3
0186a80f
01330c0f
ff66001c
149480a7
059421a7
2c0f20c6
01d30006
04542067
08942147
00060093
00d3080f
280f2026
001cfe93
0c56ff7b
00000804
08a730c3
001c0754
331cff7b
0894028c
60260093
0073640f
440f4046
08040006
0136f016
71c360c3
10f8801c
0000811c
b80c0333
680c28c3
182c8c4c
43a617c3
51b0301c
0016311c
28c34664
8c4c680c
17c306c3
301c43a6
311c51b0
46640016
c00765c3
8076e794
08040f56
0136f016
71c360c3
10f8801c
0000811c
b80c0333
680c28c3
182c8c4c
43a617c3
519c301c
0016311c
28c34664
8c4c680c
17c306c3
301c43a6
311c519c
46640016
c00765c3
8076e794
08040f56
50c33016
0404305c
10946027
10f8301c
0000311c
8c4c6c0c
155c03ac
40a614a4
518c301c
0016311c
744c4664
10946027
10f8301c
0000311c
8c4c6c0c
155c140c
40c614a4
518c301c
0016311c
355c4664
67d21831
05d2152c
14a4155c
0aa318bc
05d2154c
14a4155c
0aa318bc
05d2156c
14a4155c
0aa33ebc
05d2158c
14a4155c
0aa33ebc
1a84055c
301c0fd2
311c10f8
6c0c0000
155c8c4c
454614a4
518c301c
0016311c
055c4664
0fd21d64
10f8301c
0000311c
8c4c6c0c
14a4155c
301c4546
311c518c
46640016
08040c56
ff963016
505c40c3
005c1464
143c1444
2fc328c0
1484345c
0aa222bc
001c30c3
6007ff74
345c1a74
0ea01464
6c006017
00d36037
fff0323c
1467345c
245c1fe5
19f21464
702f6017
1444345c
700f6d00
68802017
1467345c
0c560196
00000804
40ac1016
23e464ac
23e43dd4
408c3d94
23e4648c
23e437d4
606c3794
42c3446c
30d434e4
34e442c3
604c0694
42c3444c
28d434e4
446c606c
34e442c3
604c0b94
42c3444c
069434e4
442c602c
34e442c3
606c19d4
42c3446c
169434e4
444c604c
34e442c3
602c1194
42c3442c
0c9434e4
600c4006
40c3040c
02f434e4
02c34026
00260093
00060053
08040856
01c330c3
fabc13c3
08040aa3
40c31016
ff53001c
001c8fd2
2067ff7c
301c0b35
311c10fc
6c0c0000
00066c6c
100f3664
08560006
00000804
ff967016
305c40c3
105c1464
45a21444
305c6025
001c1467
4067ff6d
01c32794
28c0143c
345c2fc3
f2bc1484
30c30aa1
ff74001c
1a746007
b0afa017
1464345c
1444245c
133cc9a2
145c0010
001c1467
ccf2ff6e
fff0353c
045c70af
48001464
6580538f
1467345c
019606c3
08040e56
008610c3
313c4306
64f2208d
5f051fe5
08041bf2
fd963016
41c300b7
6fe730c3
5f5c06b4
a40d0041
03b30026
0aa494bc
02a35006
3f5c0077
700d0021
94bc0097
203c0aa4
14c3180c
013330c3
54c38097
a0375243
00014f5c
7fe5840d
20255f05
002576f2
0c560396
00000804
460631c3
00df233c
9ebc13c3
00250aa4
00000804
408631c3
00df233c
9ebc13c3
00250aa4
00000804
462631c3
00df233c
9ebc13c3
00250aa4
00000804
fe963016
23c342c3
503c1264
a037ff00
00013f5c
00771406
03356027
00771006
53c36057
a07751a3
0f5c32c3
033c0021
04c300df
9ebc13c3
00250aa4
0c560296
00000804
7406ff96
003703a3
2f5c32c3
233c0001
01c300df
9ebc13c3
00250aa4
08040196
0208031c
031c0454
0394020c
01f30026
20d6303c
0b0d333c
fff0233c
20e6303c
0b0d333c
32a37fe5
f88c033c
00000804
019e301c
13540047
08d40047
0289301c
6b060ed2
0a940027
301c0153
008701a0
301c0654
00a7019f
60060254
080403c3
0136f016
42c351c3
219763c3
5c546007
5af42007
5854a007
56f48007
65c77408
41e45354
303c5174
6027fff0
00274db4
78082594
000626c3
049465c7
00250213
68084025
03546807
fa7401e4
071501e4
14944007
60250093
00730025
600605c3
48074008
31e40354
31e4f774
48070715
503c0594
33e30010
78089180
049465c7
b58070a0
200691a0
4cb8801c
0016811c
54a202f3
7c0c78c3
30c30d22
0001341c
440562d2
78c318a2
ec227c0c
341c37c3
62d20001
20250405
069420e4
80079fe5
0026e9d4
00060053
0f568076
00000804
0136f016
40c3fc96
62c351c3
20f72006
7f3c20b7
8f3c00c0
17c30080
35c328c3
0aa222bc
3a740007
60076097
60d73a54
207731a2
60f76025
06542027
1819365c
2f946027
04c30573
28c317c3
f2bc35c3
00070aa1
60d72374
602551a2
45d260f7
00213f5c
181d365c
25e440d7
71221a34
14946047
0010323c
51a260f7
001c4037
4027ff13
60250f94
51a260f7
182d265c
00013f5c
1825365c
001c0093
0053ff74
04960006
0f568076
00000804
0136f016
40c3fe96
82c351c3
20772006
6f3c2037
16c30040
35c32fc3
0aa222bc
76740007
16c304c3
35c32fc3
0aa222bc
6e740007
71224057
00a0331c
323c3b94
60770010
16c304c3
35c32fc3
0aa1f2bc
5e740007
71224057
00a0331c
323c2894
60770010
16c304c3
35c32fc3
0aa1f2bc
4e740007
71224057
0086331c
323c1894
60770010
16c304c3
35c32fc3
0aa1f2bc
3e740007
38c32017
16a7135c
71004057
315c18c3
60571687
00534017
6d006017
40576077
173425e4
331c7122
139400a1
0010323c
00802f3c
fe7e323c
12c304c3
35c32fc3
0aa1f2bc
1a740007
20176057
60776c80
25e44057
71221634
00a2331c
323c1294
2f3c0010
323c0080
04c3fe7e
2fc312c3
f2bc35c3
00070aa1
001c0415
0053ff74
02960006
0f568076
00000804
fe967016
51c340c3
400662c3
60094077
22946067
00803f3c
233c4026
13c3fe7e
35c32fc3
0aa1f2bc
16740007
233c6057
40770010
7fe56017
31226037
1846165c
60470006
71000b94
323c4c29
365c40ac
00061846
001c0073
0296ff74
08040e56
20c31016
10f8301c
0000311c
8c0c6c0c
12c30986
301c40e6
311c4fe0
46640016
60060dd2
602f600f
608f606f
60cf60af
616d60ef
6006614d
0856624f
00000804
60c3f016
501c71c3
511c10f8
740c0000
00ac8c4c
301c40a6
311c4fd4
46640016
8c4c740c
17c3186c
301c40c6
311c4fd4
46640016
04d218cc
3ebc17c3
18ec0aa3
17c304d2
0aa33ebc
10f8301c
0000311c
8c4c6c0c
17c306c3
301c40e6
311c4fd4
46640016
08040f56
0136f016
72c381c3
a00660c3
180c0193
824c00d3
e8bc17c3
04c30aa6
063c1bf2
a025027f
f47458e4
0f568076
00000804
0037ff96
ff53001c
13542007
46d232c3
440d5406
642d6066
40466046
602545a1
45a14026
2f5c6025
45a10001
0010033c
08040196
61c3f016
440c42c3
700f6006
64092100
16946147
0010523c
20c302a2
08350087
700c01f3
333ce429
700f43ac
20255fe5
353c59f2
6c000010
100c780f
001c0073
0f56ff74
00000804
0336f016
40c3fe96
72c391c3
440c83c3
40252122
131c4077
199400a0
00405f3c
2fc315c3
0aa1f2bc
16740007
15c304c3
38c32fc3
0aa222bc
0e740007
70802057
40177dcf
31c35def
60776d00
29c36057
0006680f
001c0073
0296ff74
0f56c076
00000804
50c33016
1f540007
0ed2014c
10f8301c
0000311c
8c4c6c0c
4646366c
4f7c301c
0016311c
158c4664
301c0ed2
311c10f8
6c0c0000
366c8c4c
301c4646
311c4f7c
46640016
08040c56
0136f016
50c3ff96
82c341c3
440c73c3
40c74122
2fc30a94
0aa1f2bc
1b740007
c017700c
700f6f00
05c3d00c
2fc314c3
22bc37c3
00070aa2
700c0e74
6d004017
2f201700
18bc28c3
700c0b25
6f00c017
0073700f
ff74001c
80760196
08040f56
40c33016
1fe651c3
29548007
20070026
524c2654
06ac4dd2
08200bd2
1f940007
0380043c
eabc268c
000708cb
04c31894
4286358c
08cbeabc
11940007
0140043c
428635ac
08cbeabc
516c0af2
652c366c
05f209a0
2085114c
08cbeabc
08040c56
ff961016
203740c3
408632c3
2f5c4c0d
4c2d0001
0020033c
401714c3
08cbb0bc
03c36017
01960045
08040856
3f36f016
a0c3f796
403771c3
7b540007
79542007
8007824c
04c37654
00601f3c
0aa4d4bc
1ac3b0c3
0080264c
00b01f3c
0aa4d4bc
40c6d0c3
00852f5c
1f3c0126
9ebc0110
903c0aa4
343c0010
3b840090
19c33d84
04c38c80
01501f3c
0aa4cabc
900080c3
1f3c04c3
cabc01a0
60c30aa4
cf3c9000
004601f0
2cc314c3
0aa50abc
700050c3
12c34017
3db431e4
1cc307c3
b0bc25c3
1e8008cb
01a01f3c
b0bc26c3
970008cb
1f3c1e00
28c30150
08cbb0bc
1e004884
01001f3c
b0bc29c3
498408cb
101c1e00
111c4f9c
41260016
08cbb0bc
1e008125
00b01f3c
b0bc2dc3
4d8408cb
1f3c1e00
2bc30060
08cbb0bc
1e004b84
03801a3c
4e4c3ac3
08cbb0bc
264c1ac3
00531080
09960006
0f56fc76
00000804
fe96f016
41c360c3
23c372c3
a1a2640c
640ca80d
640f6025
23c36809
40375d25
00013f5c
ff67201c
1cb46027
00402f3c
f2bc61d7
201c0aa1
0007ff74
a0571374
ff30353c
ff6b201c
0cb46267
500c07c3
25c33900
08cbb0bc
a057700c
700f6e80
02c34006
0f560296
00000804
0336f016
41c360c3
53c382c3
4007e1d7
00073254
60073054
640c2e54
0010233c
2cb427e4
440f61a2
2b946047
37c325c3
0aa1f2bc
25740007
4407540c
300c22b4
37e46880
00061bb4
1df420e4
07f218a2
fff0323c
700c740f
700f6025
500c08c3
540c3900
08cbb0bc
140c700c
700f6c00
01330006
ff53001c
001c00d3
0073ff7c
ff74001c
0f56c076
00000804
fe967016
503c40c3
6f3c28c0
005c0040
15c31444
345c26c3
22bc1484
00070aa2
345c2d74
706f1464
1444045c
26c315c3
1484345c
0aa222bc
20740007
245c6057
6d001464
045c708f
15c31444
0200243c
0aa2a6bc
12740007
1444345c
1484245c
03c34037
243c15c3
343c2980
fcbc2b80
30c30aa8
30e40006
001c0315
0296ff74
08040e56
fe961016
207740c3
44f202d2
ff53001c
00060553
31c32057
25b46407
280d2046
60077008
60571415
202513c3
3f5c2037
682d0001
284d2006
0030023c
405714c3
08cbb0bc
03c36057
01b30065
00211f5c
023c282d
14c30020
b0bc4057
605708cb
004503c3
08560296
00000804
0f36f016
70c3fd96
62c381c3
20b72006
4f3c2077
14c30080
00402f3c
22bc38c3
00070aa2
000bc3dc
365c6026
b4c31835
10f8901c
0000911c
60971593
433c5da2
80b70010
fff0313c
231c6077
3d940082
1bc307c3
38c32fc3
0aa1f2bc
f3dc0007
20570009
40977080
60776d20
640c19c3
01068c0c
14a4165c
301c43a6
311c4fec
46640016
000750c3
0008a2dc
680c29c3
60178c0c
0010033c
14a4165c
301c43a6
311c4fec
46640016
0007142f
60973e54
40173d80
08cbb0bc
6017542c
29a12006
540f592c
09b3b92f
0081231c
07c35294
2fc31bc3
f2bc38c3
00070aa1
40576074
20977100
60776ca0
680c29c3
01068c0c
14a4165c
301c43a6
311c4fec
46640016
000750c3
19c34c54
8c0c640c
033c6017
165c0010
43a614a4
4fec301c
0016311c
142f4664
11940007
10f8301c
0000311c
8c4c6c0c
165c05c3
43a614a4
4fec301c
0016311c
05734664
3d004097
b0bc4017
542c08cb
20066017
594c29a1
b94f540f
60574017
60776d20
6d006097
023360b7
1bc307c3
38c32fc3
0aa1f2bc
0f740007
20976017
20574c80
6d207080
40b76077
20072057
fff536dc
00730006
ff74001c
f0760396
08040f56
0136f016
40c3fe96
52c361c3
20772006
7f3c2037
17c30040
36c32fc3
0aa222bc
28740007
71224057
331c0006
24940080
0010323c
04c36077
2fc317c3
f2bc36c3
00070aa1
60571774
155c3180
40171927
1947255c
2ed0353c
06944287
b0bc03c3
000608cb
01c30133
23c312c3
0b2518bc
001c0073
0296ff74
0f568076
00000804
fe967016
61c350c3
400642c3
40374077
60876009
3f3c2494
40260080
fe7e233c
2fc313c3
f2bc36c3
30c30aa1
17746007
35004057
1967145c
245c4017
343c1987
42872d80
03c30694
08cbb0bc
01330006
12c301c3
18bc23c3
00730b25
ff74001c
0e560296
00000804
3f36f016
70c3fa96
b2c391c3
8f3ca3c3
60060180
fffc821c
680f28c3
00c0df3c
10f8c01c
0000c11c
07c30c73
2f3c18c3
39c30100
0aa222bc
5f740007
dda26157
60b76025
1f3c07c3
2dc30080
f2bc39c3
00070aa1
263c52f4
407707f0
00213f5c
04356027
00a4631c
2cc33f94
8c0c680c
1ac30206
301c43a6
311c4ffc
46640016
000750c3
2cc31d54
8c0c680c
1ac300d7
301c43a6
311c4ffc
46640016
0007142f
301c1194
311c10f8
6c0c0000
05c38c4c
43a61ac3
4ffc301c
0016311c
10664664
609703d3
40d73d80
08cbb0bc
544f40d7
00f4263c
3f5c4037
758d0001
480c2bc3
3bc3540f
6157ac0f
6d004117
61576177
9c1439e4
00730006
ff74001c
fc760696
08040f56
0f36f016
70c3fe96
52c361c3
40774006
4f3c4037
14c30040
36c32fc3
0aa222bc
2a740007
02c0a53c
0300953c
03f3b4c3
60259da2
07c36077
2fc31bc3
f2bc36c3
00070aa1
2ac319f4
00a0431c
431c0554
129400a1
605729c3
20171d80
14a4355c
0aab02bc
40176057
60776d00
36e46057
0006e014
001c0073
0296ff74
0f56f076
00000804
3f36f016
60c3f996
28f22037
3500503c
0840a03c
0480703c
503c00f3
a03c3ac0
703c1840
065c0340
365c1444
61a21464
129460c7
28c0163c
01402f3c
1484365c
0aa1f2bc
43dc0007
365c003b
21571464
365c6c80
465c1467
c63c1464
065c28c0
1cc31444
01402f3c
1484365c
0aa222bc
e3dc0007
365c0039
41571444
0e004a20
1464365c
27c32980
0b2518bc
0007d0c3
003914dc
165c6157
4c801464
60174177
202713c3
365c0b94
165c1444
6c801464
1a47365c
365c68a0
e0061a67
4f3c42b3
065c0100
1cc31444
365c24c3
46bc1484
065c0aa2
1cc31444
365c24c3
22bc1484
00070aa2
003653dc
1464365c
1444065c
602541a2
1467365c
045440c7
ff70d01c
1cc36b33
00c02f3c
1484365c
0aa1f2bc
e3dc0007
365c0034
0f3c1444
265c01a0
2d001464
b0bc4046
2f5c08cb
4aa700d1
001014dc
00d93f5c
c4dc6087
165c000f
313c1464
365c0020
265c1467
89a21444
0030313c
1467365c
607769a2
0040313c
1467365c
1cc302c3
00802f3c
1484365c
0aa1f2bc
c3dc0007
801c0031
60970000
00d0233c
0100301c
23e46fa0
801c0374
80670001
60172594
202713c3
365c0d94
265c1444
6d001464
60977baf
1f5c7bcf
165c0021
600603e5
4cf228c3
0f803ac3
4cbc101c
0016111c
b0bc4086
e08508cb
165c6026
346f1464
548f4097
808712f3
60061194
200718c3
0008c4dc
0b802ac3
4cc4101c
0016111c
b0bc24c3
e08508cb
80c70ff3
60061594
2cf218c3
0b802ac3
4ccc101c
0016111c
b0bc4066
e06508cb
165c6026
34ef1464
550f4097
80e70df3
60061594
2cf218c3
0b802ac3
4cd0101c
0016111c
b0bc4066
e06508cb
165c6026
352f1464
554f4097
81070b33
60061594
2cf218c3
0b802ac3
4cd4101c
0016111c
b0bc4086
e08508cb
165c6026
356f1464
558f4097
81470873
60061594
2cf218c3
0b802ac3
4cdc101c
0016111c
b0bc4066
e06508cb
165c6026
35af1464
55cf4097
816705b3
60061594
2cf218c3
0b802ac3
4ce0101c
0016111c
b0bc4086
e08508cb
165c6026
35ef1464
560f4097
600602f3
149480a7
28c36006
3ac34cf2
101c0f80
111c4ce8
41c60016
08cbb0bc
6026e1c5
1464165c
409734af
600754cf
000e72dc
600738c3
000e34dc
1444365c
07801ac3
1464265c
40972d00
08cbb0bc
fd806097
45471ab3
3f5c0a94
b01c00d9
80260000
0086331c
01d30c94
09944127
00d93f5c
0001b01c
331c8006
04540092
0000b01c
365c4bc3
60251464
6d0040d7
1467365c
1444065c
2f3c1cc3
365c0080
f2bc1484
00070aa1
002153dc
301c2097
4fa00100
0000901c
03f412e4
0001901c
74548007
00d0313c
047432e4
0001901c
29c301b3
3ac34bf2
101c0f80
111c4cf8
41c60016
08cbb0bc
165ce1c5
362f1464
564f4097
10f8101c
0000111c
8c0c640c
165c0106
43a614a4
517c301c
0016311c
80c34664
25540007
10f8201c
0000211c
8c0c680c
033c6097
165c0010
43a614a4
517c301c
0016311c
18c34664
0007042f
301c1394
311c10f8
6c0c0000
08c38c4c
14a4165c
301c43a6
311c517c
46640016
ff83d01c
365c3733
265c1444
2d001464
b0bc4097
38c308cb
60974c2c
29a12006
28c3794c
1951680f
24d219c3
0001901c
365c01b3
2ac31444
265c0b80
2d001464
b0bc4097
609708cb
1bc3fd80
28542007
233c6097
301c0040
6fa00100
1b1523e4
400729c3
3ac31894
101c0f80
111c4d08
40a60016
08cbb0bc
0050473c
1444365c
06001ac3
1464265c
40972d00
08cbb0bc
f1806097
1464165c
4097366f
365c568f
20971464
365c6c80
365c1467
41571464
31e412c3
ffde70dc
2ac36006
748c6ba1
0040733c
73c362f2
63d274cc
fd806085
63d2750c
fd806065
63d2754c
fd806065
63d2758c
fd806085
63d275cc
fd806065
63d2760c
fd806085
63d2764c
fd8061c5
63d2768c
fd8060a5
63d276cc
fd8061c5
10f8301c
0000311c
8c0c6c0c
0010073c
14a4165c
301c4546
311c517c
46640016
0007140f
001212dc
43c3748c
19546007
6025744c
101c744f
111c4cbc
40860016
08cbb0bc
265c740c
033c1444
746c0040
548c2980
08cbb0bc
346f2086
8c80748c
600774cc
744c1a54
744f6025
0e00740c
4cc4101c
0016111c
b0bc4086
808508cb
265c740c
0e001444
298074ac
b0bc54cc
94af08cb
908034cc
6007750c
744c1a54
744f6025
0e00740c
4ccc101c
0016111c
b0bc4066
806508cb
265c740c
0e001444
298074ec
b0bc550c
94ef08cb
9080350c
6007754c
744c1a54
744f6025
0e00740c
4cd0101c
0016111c
b0bc4066
806508cb
265c740c
0e001444
2980752c
b0bc554c
952f08cb
9080354c
6007758c
744c1a54
744f6025
0e00740c
4cd4101c
0016111c
b0bc4086
808508cb
265c740c
0e001444
2980756c
b0bc558c
956f08cb
9080358c
600775cc
744c1a54
744f6025
0e00740c
4cdc101c
0016111c
b0bc4066
806508cb
265c740c
0e001444
298075ac
b0bc55cc
95af08cb
908035cc
6007760c
744c1a54
744f6025
0e00740c
4ce0101c
0016111c
b0bc4086
808508cb
265c740c
0e001444
298075ec
b0bc560c
95ef08cb
9080360c
6007764c
744c1a54
744f6025
0e00740c
4cf8101c
0016111c
b0bc41c6
81c508cb
265c740c
0e001444
2980762c
b0bc564c
962f08cb
9080364c
6007768c
744c1a54
744f6025
0e00740c
4d08101c
0016111c
b0bc40a6
80a508cb
265c740c
0e001444
2980766c
b0bc568c
966f08cb
9080368c
600776cc
744c1a54
744f6025
0e00740c
4ce8101c
0016111c
b0bc41c6
81c508cb
265c740c
0e001444
298076ac
b0bc56cc
96af08cb
908036cc
4006740c
f42f4e21
d01c0073
0dc3ff74
fc760796
08040f56
0336f016
50c3fe96
92c361c3
4f3c83c3
20060080
fe7e143c
2fc314c3
22bc36c3
00070aa2
40574d74
60477522
323c4994
60770010
14c305c3
36c32fc3
0aa1f2bc
3e740007
54a22057
0010313c
45f26077
7fe56017
00536037
40172077
0c0c38c3
21e410c3
09c330d4
35806057
08cbb0bc
08c36017
2057600f
40774c80
60477522
323c1f94
2f3c0010
323c0080
05c3fe7e
2fc312c3
f2bc36c3
00070aa1
40171174
0c0c6297
21e410c3
02570ed4
35806057
08cbb0bc
02972017
0006200f
001c00d3
0073ff74
ff7c001c
c0760296
08040f56
0136f016
60c3fc96
43c351c3
826482c3
ff53201c
6c540007
b8bc2a06
9a6f0b06
5254a007
153c06c3
42860480
08cbb0bc
0140063c
05c0153c
b0bc4286
701c08cb
711c10f8
7c0c0000
055c8c0c
3a6c15c4
301c4646
311c4f8c
46640016
5066194f
46540007
2980153c
15c4255c
08cbb0bc
15c4355c
055c796f
00071664
355c2554
60071644
7c0c2154
3a6c8c0c
301c4646
311c4f8c
46640016
0df2198f
8c4c7c0c
3a6c194c
301c4586
311c4f8c
46640016
03d35066
1644155c
1664255c
08cbb0bc
1664355c
38c379af
11546007
16bc0fc3
0df20b1c
163c0fc3
42060380
0b1bf6bc
620603f2
0fc37a4f
0b1c08bc
02c34006
80760496
08040f56
40c3f016
62c351c3
01c373c3
4f062006
0891b0bc
200604c3
b0bc4c06
7fe60891
b26f700f
f2efd2cf
08040f56
70c3f016
52c341c3
426463c3
200602c3
b0bc4486
82e70891
1c090e94
0aa1d0bc
05350087
076c301c
039374af
07d0201c
031354af
1da2780c
0aa1d0bc
3e87303c
6d0054ac
780c74af
780f6025
d0bc1da2
303c0aa1
54ac0647
74af6d00
6025780c
053c780f
17c30140
d6bc26c3
74ac0aa1
f894321c
053c74af
17c30100
d6bc26c3
748c0aa1
748f7fe5
00c0053c
26c317c3
0aa1d6bc
0080053c
26c317c3
0aa1d6bc
0040053c
26c317c3
0aa1d6bc
17c305c3
d6bc26c3
00260aa1
08040f56
40c31016
100f0006
104f102f
138f110f
13cf13af
045c0186
000603e5
0407045c
1835045c
112f0006
116f114f
045c118f
045c0425
145c0c25
20061447
1467145c
1487245c
14a7345c
2980043c
b0bc4406
60060891
15c7345c
15e7345c
1607345c
1627345c
1647345c
1667345c
1687345c
16a7345c
2d80043c
42862006
0891b0bc
045c0006
043c1765
20062ed0
b0bc4286
20060891
180d145c
183d145c
345c6006
145c1846
145c1855
145c185d
145c181d
145c1825
2006182d
19c7145c
19e7145c
1a07145c
1a27145c
3500043c
b0bc4b86
043c0891
20063ac0
b0bc4b86
60060891
1865345c
186d345c
1875345c
187d345c
1885345c
1895345c
189d345c
18a5345c
045c0006
045c18c7
045c18e7
045c1907
045c1927
045c1947
045c1967
345c1987
045c1815
085619a7
00000804
3f3cff96
40060040
fe7e233c
2fc312c3
0ace82bc
03740007
63f26017
ff7b001c
08040196
3f36f016
70c3fd96
d2c351c3
000793c3
001092dc
62dc2007
40070010
001032dc
02dc6007
2f3c0010
22bc0040
00070aa2
000fc3dc
15c307c3
00802f3c
0aa26abc
33dc0007
740c000f
60255da2
4087740f
40c70654
40e70454
000e84dc
0040cf3c
15c307c3
39c32cc3
0aa1f2bc
d3dc0007
601c000d
6057ff7c
96dc6847
801c000d
811c10f8
18c30000
8c0c640c
20060866
301c44c6
311c4fbc
46640016
d066b0c3
52dc0007
28c3000c
8c0c680c
0086001c
44c62006
4fbc301c
0016311c
a0c34664
18c30ef2
8c4c640c
1ac30bc3
301c44c6
311c4fbc
46640016
1533d066
00248f5c
540c0bc3
28c33d00
08cbb0bc
2057740c
540f4c80
331c7d22
2f9400a0
0010323c
07c3740f
2cc315c3
f2bc39c3
00070aa1
740c6e74
60255da2
601c740f
40c7ff70
07c36894
2cc315c3
f2bc39c3
30c30aa1
30e40006
0b730715
5da2740c
60250100
4057740f
fff0323c
57f26077
0ab192bc
ff54601c
4d740007
5da2740c
740f6025
ff55601c
00a1231c
4f3c4494
07c30040
24c315c3
f2bc39c3
00070aa1
740c3874
60255da2
601c740f
4067ff6d
07c33294
24c315c3
f2bc39c3
00070aa1
20572874
ff66601c
25f42007
5da2740c
740f6025
ff6e601c
1d944007
fff0413c
ff7c601c
0085431c
0ac316d4
24c33d80
08cbb0bc
4057740c
740f6d00
0007df5c
18c30bc3
34c32ac3
0ad04abc
007360c3
ff74601c
10f8501c
0000511c
8c4c740c
20060bc3
301c44c6
311c4fbc
46640016
8c4c740c
20060ac3
301c44c6
311c4fbc
46640016
601c00d3
0073ff53
ff74601c
039606c3
0f56fc76
00000804
ff963016
42c330c3
a037a006
20a7a80f
0010b2dc
13b420a7
f2dc2047
2047000c
200707b4
20272254
001c94dc
20670ad3
000e12dc
24dc2087
1c13001c
12dc2107
21070018
20c708b4
000ff2dc
64dc20e7
2d13001b
42dc2147
21470018
0017a0dc
c4dc2167
3413001a
019f031c
031c2c54
08b4019f
1b540b07
019e031c
0019f4dc
031c03b3
09540286
0289031c
031c0b54
44dc01a0
03930019
5018301c
0016311c
201c1073
211c5020
2f730016
5028501c
0016511c
40a6a037
301c16b3
311c5030
0c330016
503c201c
0016211c
501c2e93
511c5048
0a130016
0286031c
031c3554
17b40286
020c031c
031c5654
09b4020c
0205031c
031c2454
04dc0208
08d30016
020d031c
031c4d54
84dc020e
0a130015
028f031c
031c2854
09b4028f
0288031c
031c1854
a4dc0289
03130014
0290031c
031c1f54
24dc0291
04330014
5054301c
0016311c
201c0a93
211c505c
26730016
5068501c
0016511c
301c01f3
311c5074
02330016
5080201c
0016211c
501c2493
511c508c
a0370016
0a934126
5098301c
0016311c
a1266037
201c0233
211c50a4
04330016
50ac501c
0016511c
301c0833
311c50b4
60370016
b00fa106
201c20f3
211c50bc
1eb30016
0206031c
031c1454
0c540285
0203031c
000f94dc
50c4201c
0016211c
60e64037
501c1e13
511c50cc
f9530016
50d8301c
0016311c
a0e66037
1fc3fbb3
0ace82bc
08a71c33
031c0654
c4dc028c
0113000d
50e0201c
0016211c
60a64037
501c1a53
511c50e8
a0370016
500f4106
0ea71973
0ec70554
000c74dc
301c00d3
311c50f0
f4b30016
50fc201c
0016211c
031c1713
65540090
0090031c
031c16b4
4c540081
0081031c
08a708b4
031c3354
a4dc0080
0713000a
0083031c
031c2154
24dc0085
02f3000a
0095031c
031c2854
09b40095
0091031c
031c1854
44dc0092
04f30009
0097031c
031c3554
c4dc00a8
05330008
5108301c
0016311c
201c05f3
211c510c
06330016
5110501c
0016511c
301c03d3
311c5114
ed930016
511c201c
0016211c
501c0453
511c5120
01f30016
5124301c
0016311c
201c0233
211c5128
02730016
512c501c
0016511c
4066a037
301cf1f3
311c5130
60370016
e993a066
5134201c
0016211c
60664037
0e870993
0ea70454
00d34994
5138301c
0016311c
201ce733
211c5140
06330016
0092031c
201c3b94
211c5148
03130016
349409e7
514c201c
0016211c
09070453
09071754
08e704b4
01b31f94
155409e7
0097031c
201c1994
211c5154
40370016
03736086
5158501c
0016511c
301ce933
311c5160
e1130016
5168201c
0016211c
61064037
331c0153
08940294
5170201c
0016211c
61264037
0017700f
0c560196
00000804
0f36f016
50c3fc96
42c391c3
4ed2a3c3
04944027
0aa51abc
804709d2
531c0494
04540285
0000801c
801c0073
3f3c0002
20060100
fe7e133c
14c305c3
c0bc23c3
70c30ab2
3854e007
0080bf3c
1bc300d7
0aa49ebc
2ac360c3
688020d7
38846025
00204f3c
14c30c00
0aa4cabc
502140c6
0010503c
14c309c3
b0bc25c3
39c308cb
1bc30e80
b0bc26c3
b70008cb
868019c3
17c304c3
b0bc40d7
28c308cb
20d749d2
40a67080
20d74c0d
40067080
18c34c2d
650040d7
04960e80
0f56f076
00000804
3f36f016
40c3b296
407791c3
1f3c0b06
40061240
a2bc32c3
d0c30ab4
228604c3
05102f3c
0aa828bc
043cc0c3
22860140
00802f3c
0aa828bc
114cb0c3
2f3c316c
84bc0d40
a0c30aa9
83c3724c
04c368d2
09a01f3c
3ebc44a6
80c30aa8
3d843cc3
2ac33b84
6f3cad00
808610b0
11007f3c
16c305c3
0aa4cabc
4b9d073c
8047b400
58840294
df659fe5
f3949fe7
ff7c001c
23c36057
42b452e4
11006f3c
0f707f3c
2f3ca006
40371240
024f463c
0e8039c3
24c317c3
08cbb0bc
e0a5b600
32c34017
f39463e4
0a8029c3
2dc316c3
08cbb0bc
95803dc3
0a0029c3
05101f3c
b0bc2cc3
4c8408cb
0e0039c3
00801f3c
b0bc2bc3
4b8408cb
0a0029c3
0d401f3c
b0bc2ac3
4a8408cb
69d238c3
0a0029c3
09a01f3c
b0bc28c3
488408cb
4e9604c3
0f56fc76
00000804
0f36f016
70c3e796
bf3c43c3
01c30020
2bc312c3
0aa828bc
8f3ca0c3
04c304b0
400618c3
a2bc32c3
50c30ab4
9a8490c3
05f06f3c
16c309c3
0aa4cabc
07c340c3
24c316c3
08cbb0bc
18c31e00
b0bc25c3
728008cb
1bc31d80
b0bc2ac3
39c308cb
19960e00
0f56f076
00000804
0336f016
60c3fd96
52c371c3
240c83c3
40062077
60a2540f
ff70201c
409460c7
0010313c
00c02f3c
fc7e323c
2f3c12c3
62970080
0aa1f2bc
ff74201c
30740007
00249f5c
80078097
f90c343c
7f526e20
01134383
58a2740c
740f6d00
0010313c
40976077
fff0323c
205760b7
3c0f54f2
000c831c
140c1454
2fc318c3
0ab2c0bc
0dd210c3
34e46017
39c30794
24c31980
08cbeabc
201c04d2
0053ff6c
02c34006
c0760396
08040f56
0f36f016
50c3fc96
82c391c3
240c73c3
40a220f7
00a1231c
213c6a94
4f3c0010
243c0100
6f3cfe7e
14c30080
f2bc26c3
00070aa1
05c35c74
26c314c3
22bc37c3
00070aa2
60975474
20d7a3c3
bf3ca184
08d30040
14c305c3
37c326c3
0aa222bc
45740007
60776006
05c3e037
2bc314c3
cabc60a6
00070ab5
40d73a74
60277522
323c0494
60f70030
752240d7
2f946087
0010323c
05c360f7
26c314c3
f2bc37c3
00070aa1
60572474
16946ec7
752240d7
1d946087
0010323c
05c360f7
26c314c3
f2bc37c3
00070aa1
20d71274
28c37480
60976a8f
60d76aaf
6c802097
60d760f7
b9143ae4
700f49c3
00730006
ff74001c
f0760496
08040f56
0736f016
50c3fc96
92c341c3
40f74006
6f3c40b7
7f3c00c0
16c30080
34c327c3
0aa222bc
36150007
05c307b3
27c318c3
22bc34c3
00070aa2
60063574
80376077
18c305c3
60e62ac3
0ab5cabc
2a740007
d5a260d7
60f76025
18c305c3
34c327c3
0aa1f2bc
1e740007
0086631c
60570e94
0b946e87
39c34097
1667235c
750040d7
325c29c3
01931647
409760d7
60f76d00
86c30093
0040af3c
34e460d7
0006c714
001c0073
0496ff74
0f56e076
00000804
0136f016
70c3f896
42c361c3
02005f3c
253c4006
15c3fe7e
01402f3c
22bc36c3
00070aa2
41d74974
345c7d00
615718c7
18e7345c
5f3c85c3
07330180
07c3c037
25c318c3
cabc6146
00070ab5
61973574
19546907
04b46907
249468e7
69e701b3
331c1954
1e940097
1859345c
61376372
00812f5c
345c02b3
60721859
2f5c60f7
01d30061
1859345c
60b76172
00412f5c
345c00f3
62721859
2f5c6077
245c0021
345c185d
60251904
1907345c
36e461d7
0006c614
001c0073
0896ff74
0f568076
00000804
1f36f016
50c3fa96
21772006
1604805c
15e4605c
28c3c3d2
001c44f2
2413ff53
331c7809
a4dc00a3
4f3c0011
40260180
fe7e243c
01007f3c
14c306c3
38c327c3
0aa1f2bc
a3dc0007
06c30010
27c314c3
22bc38c3
00070aa2
001013dc
0000901c
bf3ca4c3
cf3c00c0
1dd30080
1ac306c3
38c327c3
0aa222bc
03dc0007
4006000f
8f5c40f7
06c30007
2bc31ac3
cabc60c6
00070ab5
000e53dc
99a26157
14948027
40b74006
61776025
1ac306c3
38c32cc3
0aa1f2bc
23dc0007
6157000d
602559a2
80776177
400643f2
41574077
60877922
000c54dc
0010323c
06c36177
27c31ac3
f2bc38c3
00070aa1
000b93dc
331c60d7
22dc0090
331c0009
16b40090
0081331c
331c6d54
08b40081
375468a7
0080331c
000934dc
331c0ab3
36540083
0085331c
0008b4dc
331c02b3
3c540095
0095331c
331c08b4
1a540091
0092331c
10137d94
0097331c
331c5954
769400a8
60260f33
1865355c
00211f5c
186d155c
19004157
25c32117
0aa5b2bc
41570c93
21171900
08bc25c3
0bb30aa6
19004157
25c32117
0ab69abc
40260ad3
1875255c
00213f5c
187d355c
18802157
25c32117
0aa9babc
60260713
180d355c
00211f5c
1885155c
19004157
25c32117
0aaa8ebc
40260753
1765255c
00213f5c
1895355c
18802157
25c32117
0aaacebc
60260393
183d355c
00211f5c
189d155c
19004157
25c32117
0aa698bc
402603d3
1855255c
00213f5c
18a5355c
18802157
25c32117
0ab6f2bc
16150007
60260473
1815355c
00211f5c
188d155c
19004157
25c32117
0aab84bc
06150007
40570273
901c43d2
61570001
6c802117
61576177
10dc38e4
001cfff1
39c3ff60
09c365f2
001c0073
0696ff74
0f56f876
00000804
0336f016
50c3fd96
62c391c3
e29783c3
00c04f3c
143c240c
4006fc7e
14c3580f
00802f3c
22bc37c3
30c30aa2
ff74001c
1e746007
05c3e037
26c314c3
cabc38c3
30c30ab5
ff70001c
12746007
75224057
0a9460a7
0010323c
001c6077
55a2ff6e
602547f2
20576077
2c0f39c3
03960006
0f56c076
00000804
fb96f016
61c350c3
01404f3c
143c2006
7f3cfe7e
14c30040
36c327c3
0aa222bc
41740007
14c305c3
00802f3c
0aa26abc
39740007
05c3c037
2f3c14c3
604600c0
0ab888bc
2f740007
75224117
109460c7
0010323c
05c36137
27c314c3
f2bc36c3
00070aa1
61172074
6c802057
41176137
60877522
323c1894
2f3c0010
323c0140
05c3fe7e
2f3c12c3
36c30040
0aa1f2bc
09740007
611705c3
40573580
08cbb0bc
00730057
ff74001c
0f560596
00000804
fe967016
403c50c3
6f3c28c0
005c0040
14c31444
355c26c3
22bc1484
00070aa2
000993dc
1444355c
1484255c
03c34037
253c14c3
604601c0
0ab888bc
a3dc0007
74ec0008
0206331c
201c2954
331cff6c
84dc0285
355c0008
055c1464
41a21444
355c6025
40671467
14c37894
355c26c3
f2bc1484
00070aa1
255c6d74
355c1464
2d221444
0010323c
1467355c
68942007
cabc05c3
20c30aa3
355c0cb3
255c1444
40371484
14c303c3
3340253c
cabc6066
00070ab5
055c4f74
92bc19a4
201c0ab1
0007ff54
355c4f74
055c1464
41a21444
355c6025
40671467
14c34094
355c26c3
f2bc1484
00070aa1
355c3574
255c1464
c9a21444
355c6025
c0071467
60573194
fff0233c
301c4077
311c10f8
6c0c0000
02c38c0c
14a4155c
301c40c6
311c5184
46640016
5066140f
1c540007
1444355c
1464255c
40572d00
08cbb0bc
744f6026
342f2057
1464355c
355c6c80
26c31467
201c0133
00d3ff74
ff6d201c
201c0073
02c3ff6e
0e560296
00000804
3f36f016
50c3fe96
62c32037
02c383c3
0af286bc
08c390c3
0af286bc
06c3c0c3
0ae318bc
08c3b0c3
0ae318bc
7bc3d0c3
a0c37984
4ac3ac84
033c7380
233c0040
20170060
101c640c
2077ff53
341432e4
cabc15c3
20460aa4
403c3421
07c30010
9ebc3600
90000aa4
44d229c3
76216006
06c38025
60bc3600
00770af2
1c940007
70801bc3
55a14046
0010433c
36000ac3
0aa49ebc
3cc38200
1f5c65d2
36210021
08c38025
60bc3600
00770af2
2dc305f2
80177100
0057700f
fc760296
08040f56
3f36f016
80c3fe96
000791c3
000c02dc
d2dc2007
c0ec000b
4b54c007
60477989
29c31a94
0293e92c
04c39c2c
08920ebc
336430c3
384cb82c
00462037
23c314c3
4abc35c3
00070aa5
000a24dc
e007fc0c
05b3ec94
1a946027
ed4c39c3
9c2c0293
0ebc04c3
30c30892
b82c3364
2037384c
14c30026
35c323c3
0aa54abc
74dc0007
fc0c0008
ec94e007
60870253
39c31094
1a64235c
31c3384c
099423e4
015c19c3
382c1a44
08cbeabc
71540007
f6b3d80c
e8cc28c3
e0070026
801c6b54
c8c30000
00278f5c
a8c3b8c3
7d89d8c3
1c946047
c92c29c3
1554c007
0001801c
982c0253
0ebc04c3
30c30892
bc2c3364
20373c4c
14c30046
35c323c3
0aa54abc
d80cc0c3
ee94c007
60270673
19c31b94
c007c54c
60771454
982c0253
0ebc04c3
30c30892
bc2c3364
40375c4c
14c30046
35c323c3
0aa54abc
d80cb0c3
ee94c007
608702f3
29c31594
1a44025c
225c0fd2
7c4c1a64
21e413c3
3c2c0994
08cbeabc
a01c05f2
dac30001
a01c0073
fc0c0001
ae94e007
43d228c3
6bd23cc3
23d22057
47d22bc3
00163d3c
0a3ca383
00530016
02960006
0f56fc76
00000804
e996f016
72c360c3
20371264
05770006
04f70537
10fc301c
0000311c
6c6c6c0c
05b73664
2f5c06c3
12c30001
02802f3c
05403f3c
0ab09ebc
92dc0007
2557000c
323c58a2
7fe502b6
63f27f32
1f9445a7
53c37fe5
313ca072
65770010
05404f3c
05000f3c
24c316c3
0aa1d6bc
04c00f3c
24c316c3
0aa1d6bc
333c6517
24d703c7
333c6c80
233c03c7
00b3528d
f4dc4b47
23c30009
6d206597
6f3c65b7
06c30040
9cbc2486
501c08cb
511c10fc
740c0000
0f3c6c8c
36640580
0bb4301c
0000311c
8e2c6c2c
78127209
111c2006
31831000
67546007
6c0c740c
0aa9035c
035c10c3
203c0ab1
135c40ac
213c0ab9
035c812c
203c0ac1
4077c12c
0ac9135c
135c01c3
213c0ad1
035c402c
203c0ad9
135c812c
213c0ae1
40b7c12c
0ae9035c
035c10c3
203c0af1
135c40ac
213c0af9
035c812c
203c0b01
40f7c12c
0b09135c
135c01c3
213c0b11
035c402c
203c0b19
135c812c
213c0b21
4137c12c
0b29035c
035c10c3
203c0b31
135c40ac
213c0b39
035c812c
203c0b41
4177c12c
0b49135c
135c01c3
213c0b51
035c402c
203c0b59
135c812c
313c0b61
321cc12c
61b7f894
007306c3
15540007
02801f3c
40bce8f2
00070aa4
52091054
00d332c3
0aa3fabc
12090ad2
361c30c3
033c0010
0093090b
00530006
17960026
08040f56
0f36f016
40c3fb96
82c3b1c3
5f3c73c3
240c0140
fe7e153c
15c3ca6c
00402f3c
0aa222bc
03dc0007
af5c000f
9f3c0084
04c30080
29c315c3
22bc37c3
30c30aa2
23dc6007
04c3000e
29c315c3
22bc37c3
00070aa2
000d93dc
04c3e037
2f3c15c3
618600c0
0ab888bc
e3dc0007
4117000c
60877122
000c94dc
0010323c
04c36137
29c315c3
f2bc37c3
00070aa1
000bd3dc
71004117
618f08c3
21176097
41374c80
60877122
000b14dc
0010323c
04c36137
29c315c3
f2bc37c3
00070aa1
000a53dc
71004117
61af08c3
20976117
61376c80
04c3e037
263c15c3
363c0040
fcbc0240
00070aa8
000913dc
51a26117
61376025
0082231c
231c1b54
075400a1
0080231c
000834dc
02734006
794f6026
1f3c04c3
2f3c0100
37c30080
0aa1f2bc
600730c3
61177374
6c802097
404600b3
6117594f
61376025
02c0563c
01008f3c
04c3e037
25c318c3
06c0363c
0aa8c6bc
600730c3
05c35b74
0361165c
febc4006
301c0aba
0007ff6a
41175354
68a01ac3
10c30057
271531e4
331c7122
239400a0
0010323c
04c36137
2f3c18c3
37c30080
0aa1f2bc
3a740007
04c0563c
04c3e037
25c318c3
06d0363c
0aa8c6bc
2e740007
165c05c3
40260369
0abafebc
ff69301c
26540007
0ac34117
20576820
30e401c3
71221815
00a1331c
323c1494
2f3c0010
323c0140
04c3fe7e
2f3c12c3
37c30080
0aa1f2bc
0a740007
00976117
61376c00
1bc34117
6006440f
301c0073
03c3ff74
f0760596
08040f56
0336f016
50c3fc96
62c391c3
e40c83c3
01004f3c
fe7e743c
582f4380
2f3c14c3
22bc0080
00070aa2
60975974
40d76fa0
784f6d00
331c7522
0d9400a0
0020323c
05c360f7
2f3c14c3
6abc0040
00070aa2
08930415
60776006
352240d7
321c31c3
6027ff5f
323c3bb4
4f3c0010
343c0100
05c3fe7e
2f3c14c3
38c30080
0aa1f2bc
2c740007
209760d7
60f76c80
00078f5c
14c305c3
00c0263c
02c0363c
0aa8c6bc
1c740007
14c305c3
38c326c3
0abbeabc
14740007
6fa060d7
12c3584c
093431e4
14c305c3
38c326c3
0ab61ebc
06740007
39c320d7
00062c0f
001c0073
0496ff74
0f56c076
00000804
f596f016
61c340c3
1444305c
005c27f2
6c001464
19c7345c
205c00d3
6d001464
1a07305c
1464545c
1444045c
607762a2
0010353c
1467345c
27c3e057
40375d25
00013f5c
ff67101c
3bb46027
28c0143c
02802f3c
1484345c
0aa1f2bc
101c30c3
6007ff74
42972e74
ff30323c
ff6b101c
27b46267
1444345c
00800f3c
1464745c
b0bc2f80
629708cb
1464045c
345c6c00
6ea01467
345cc4f2
007319e7
1a27345c
00800f3c
00212f5c
26c312c3
0abafebc
07f22006
0b0d363c
7f327fe5
f690133c
0b9601c3
08040f56
ff967016
61c350c3
1444005c
28c0153c
355c2fc3
22bc1484
401c0aa2
0007ff74
05c31474
68bc2006
00070abd
401c0415
c2f2ff6a
05c38006
68bc2026
00070abd
c3d20415
ff69401c
019604c3
08040e56
ff963016
51c340c3
0aa942bc
2f740007
1444345c
1484245c
03c34037
28c0143c
0180243c
88bc6026
00070ab8
04c32074
c6bc2006
00070aab
04c31a74
ccbc15c3
50c30abd
202604c3
0aabc6bc
0f740007
1cbc04c3
00070ab9
353c0a74
25c3fff0
32c323a3
53837f52
05c3a2d2
0c560196
00000804
0136f016
71c340c3
83c362c3
0007a197
40073154
a0072f54
60062d54
0407355c
5ebc05c3
52460ae2
26940007
14c305c3
e8bc27c3
03d20ae4
02f305c3
0100453c
5ebc04c3
06d20ae2
7ebc05c3
52460ae2
04c30273
28c316c3
0ae4e8bc
0cd220c3
7ebc05c3
04c30ae2
0ae27ebc
ff72201c
201c0073
02c3ff53
0f568076
00000804
fe967016
42c351c3
4c0c63c3
71224077
36946047
0010323c
00802f3c
fe7e323c
12c304c3
61972fc3
0aa1f2bc
28740007
00070017
20570cf4
313c50a2
60770010
303c45f2
6037fff0
20770053
5ebc05c3
72460ae2
16940007
405705c3
40173100
0ae4e8bc
05c307d2
0ae27ebc
ff72301c
60170133
6c802057
30c3780f
301c0073
03c3ff74
0e560296
00000804
fd96f016
61c350c3
73c342c3
00402f3c
0aa222bc
5e740007
16c305c3
00802f3c
0aa26abc
56740007
345c6026
e0370407
14c304c3
36c325c3
0abe6ebc
4d740007
04c3e037
0100143c
36c325c3
0abe6ebc
43740007
04c3e037
0200143c
36c325c3
0abe6ebc
39740007
04c3e037
0300143c
36c325c3
0abe6ebc
2f740007
04c3e037
0400143c
36c325c3
0abe6ebc
25740007
04c3e037
0500143c
36c325c3
0abe6ebc
1b740007
04c3e037
0600143c
36c325c3
0abe6ebc
11740007
04c3e037
0700143c
36c325c3
0abe6ebc
000630c3
071530e4
001c0093
0073ff74
ff71001c
0f560396
00000804
fe967016
41c350c3
280c62c3
50a22077
31944047
0010213c
00801f3c
fe7e213c
2fc304c3
0aa1f2bc
25740007
50a22057
0010313c
45f26077
7fe56017
00536037
05c32077
0ae25ebc
00077246
05c31694
31806057
e8bc4017
07d20ae4
7ebc05c3
301c0ae2
0133ff72
40576017
780f6d00
007330c3
ff74301c
029603c3
08040e56
0136f016
70c3fe96
62c341c3
200683c3
20372077
00405f3c
2fc315c3
22bc34c3
00070aa2
60571874
601751a0
13b432e4
17c306c3
34c325c3
0abf26bc
0b740007
17c308c3
34c325c3
0abf26bc
000630c3
031530e4
ff55001c
80760296
08040f56
fe96f016
51c340c3
73c362c3
00402f3c
0aa222bc
38740007
15c304c3
6abc2fc3
00070aa2
06c33174
25c314c3
26bc37c3
00070abf
063c2c74
14c30100
37c325c3
0abf26bc
23740007
0200063c
25c314c3
26bc37c3
00070abf
063c1a74
14c30300
37c325c3
0abf26bc
11740007
0400063c
25c314c3
26bc37c3
00070abf
60260874
00067a8f
001c00d3
0073ff74
ff62001c
0f560296
00000804
ff96f016
71c360c3
53c342c3
22bc2fc3
30c30aa2
ff74001c
2a746007
16c304c3
35c327c3
0abf26bc
20740007
0100043c
27c316c3
26bc35c3
00070abf
043c1774
16c30200
35c327c3
0abf26bc
0e740007
0300043c
27c316c3
26bc35c3
00070abf
60060574
03c3728f
001c0073
0196ff62
08040f56
ff96f016
71c360c3
53c342c3
22bc2fc3
30c30aa2
ff74001c
16746007
16c304c3
35c327c3
0abf26bc
0c740007
0100043c
27c316c3
26bc35c3
30c30abf
30e40006
001c0315
0196ff62
08040f56
0136f016
50c3ff96
82c341c3
2fc363c3
0aa222bc
600730c3
60065e74
325c28c3
700c0407
604775a2
05c34154
2fc314c3
22bc36c3
00070aa2
05c34e74
26c314c3
0aa2b8bc
600730c3
500c4674
123c7522
300f0010
099460a7
313c54a2
700f0010
ff6e001c
079343d2
700c500f
602555a2
001c700f
4067ff6d
05c33394
2fc314c3
f2bc36c3
30c30aa1
25746007
54a2300c
0010313c
42d2700f
05c3300f
2fc314c3
22bc36c3
00070aa2
08c31674
24c315c3
26bc36c3
30c30abf
10746007
0100083c
24c315c3
26bc36c3
30c30abf
30e40006
00930715
ff74001c
001c0073
0196ff71
0f568076
00000804
3f36f016
70c3fa96
40f781c3
9f5c60b7
df5c0224
a5170264
10f8301c
0000311c
8c0c6c0c
20060806
301c44c6
311c4fa8
46640016
60c3b0c3
d2dc0007
531c0017
4754020e
020e531c
531c12b4
2d540208
0208531c
531c05b4
51940205
531c04d3
2d54020c
020d531c
07b34a94
028f531c
531c2654
08b4028f
0288531c
531c0c54
3d940289
531c0253
2d540290
0291531c
03f33694
18c307c3
d2bc2bc3
a01c0b05
c01c0289
05130010
18c307c3
18bc2bc3
a01c0b25
c01c0058
03d30014
18c307c3
c6bc2bc3
a01c0b24
c01c019e
02930020
18c307c3
6ebc2bc3
a01c0b24
c01c01a0
01530040
18c307c3
16bc2bc3
a01c0b24
c01c019f
00070030
001162dc
10f8301c
0000311c
8c4c6c0c
20060bc3
301c44c6
311c4fa8
46640016
21b3c006
61776006
10f8401c
0000411c
ac0c700c
0098001c
44c62006
4fa8301c
0016311c
70c35664
ac0c700c
0200001c
44c62006
4fa8301c
0016311c
80c35664
8c0c700c
0200001c
44c62006
4fa8301c
0016311c
90c34664
28c3e5d2
000743d2
efd23394
10f8301c
0000311c
8c4c6c0c
200607c3
301c44c6
311c4fa8
46640016
6fd238c3
10f8301c
0000311c
8c4c6c0c
200608c3
301c44c6
311c4fa8
46640016
400729c3
000a42dc
10f8301c
0000311c
8c4c6c0c
200609c3
301c44c6
311c4fa8
46640016
07c31293
f4bc2557
00070b1c
d31c2f94
2cb40200
1f3c00d7
27c30140
42bc6097
00070ac0
08c32374
2dc32497
08cbb0bc
1dc308c3
01002f3c
72bc37c3
60c30b1c
a2dc1287
00070008
09c31274
2cc31bc3
94bc3ac3
06e40ab5
01170a94
26c319c3
08cbeabc
c02604f2
c0060053
e6bc07c3
401c0b1c
411c10f8
700c0000
07c3ac4c
44c62006
4fa8301c
0016311c
700c5664
08c3ac4c
44c62006
4fa8301c
0016311c
700c5664
09c38c4c
60060713
301c6137
311c10f8
6c0c0000
0a068c0c
44c62006
4fa8301c
0016311c
50c34664
2d540007
0ace6cbc
29740007
209700d7
46bc25c3
00070ad0
3f3c0f74
60370100
0497a077
2bc31dc3
f4bc3cc3
04f20ade
c027c117
c0060254
b6bc05c3
301c0ad2
311c10f8
6c0c0000
05c38c4c
44c62006
4fa8301c
0016311c
00534664
301cc006
311c10f8
6c0c0000
0bc38c4c
44c62006
4fa8301c
0016311c
01334664
0206931c
931caf54
eb940285
0013ded3
069606c3
0f56fc76
00000804
0736f016
60c3fa96
42c351c3
12c393c3
0abdf4bc
a01c20c3
2ae40000
323c0715
60270970
000c05dc
165ca2c3
801c1464
588c0000
13e432c3
790c2434
ff73201c
17dc6027
365c000b
6c801444
15e7365c
265c788c
6d201464
1607365c
1627165c
54bc06c3
20c30ab7
0000801c
061508e4
ff60231c
000984dc
388c82c3
1467165c
1444365c
1484265c
03c34037
28c0163c
01402f3c
88bc6026
20c30ab8
33dc0007
06c30008
0aa45cbc
400720c3
201c7c74
6157ff68
01c338cc
759430e4
1761165c
180c2cf2
382c0ad2
263c28d2
18bc2d80
20c30b25
67940007
5f548007
5d54a087
5b54a1c7
1809065c
301c0ed2
311c10f8
6c0c0000
09c36cac
2ed0163c
70c33664
10940007
10fc301c
0000311c
6d4c6c0c
163c09c3
36640480
201c70c3
0007ff44
165c4254
2dd21819
4bd25d69
40075d49
365c3854
65d21821
1829365c
313432e4
3c0c1c6c
05c0263c
0b2518bc
000720c3
80272a94
786c2294
1444265c
9c6c388c
1c2cbc0c
1b8c0037
18ac0077
18cc00b7
065c00f7
013714a4
25a00980
35c324c3
0ac0b6bc
ff65201c
07c30ed2
32bc16c3
201c0aba
07d2ff3a
45f22ac3
007328c3
ff12201c
069602c3
0f56e076
00000804
50c37016
0ac256bc
000760c3
17cc4474
1ef40007
10f8301c
0000311c
8c0c6c0c
155c0025
40a614a4
500c301c
0016311c
40c34664
2e540007
57cc37ac
08cbb0bc
400677cc
97af51a1
355c6026
74ec0407
0285331c
740c2094
1d546007
0007142c
301c1a54
311c10f8
6c0c0000
155c8c0c
40c614a4
500c301c
0016311c
40c34664
340c09d2
b0bc542c
940f08cb
744f6026
d0660053
0e5606c3
00000804
0736f016
fbd8f21c
91c350c3
73c362c3
2244af5c
42804f3c
143c240c
14c3fc7e
42402f3c
0aa222bc
93dc0007
3f5c0009
83c32124
21041f5c
001c8184
87e4ff66
000935dc
14c305c3
37c326c3
0abcf4bc
53dc0007
e0370008
14c305c3
0480263c
88bc6026
00070ab8
3f5c7a74
55a22104
3f5c6025
40672107
3f3c1a94
20064280
fa7e133c
14c305c3
37c323c3
0aa1f2bc
65740007
20e43f5c
1f5c7a2f
74802104
2f5c7a0f
650020e4
21073f5c
21043f5c
343438e4
1f3c05c3
26c34200
72bc37c3
00070aa7
5f3c4c74
05c30140
59ec39cc
22643f5c
0ab0fcbc
200605c3
3ac34026
0ac256bc
40740007
584c782c
20372317
20773a0c
20b73a2c
20f73a4c
21372006
12c303c3
61974157
0ac0b6bc
05c340c3
0aa364bc
1d948007
0ac304b3
0ebc39ac
00070ba7
782c1f54
806c584c
202ca00c
3a0c2037
3a2c2077
3a4c20b7
200620f7
03c32137
24c312c3
b6bc35c3
0ad20ac0
21043f5c
680f29c3
00d30006
ff74001c
001c0073
f21cff41
e0760428
08040f56
0736f016
70c3fb96
a2c391c3
21372006
01404f3c
fc7e143c
c2eca2cc
01008f3c
14c305c3
36c328c3
0aa222bc
53740007
14c305c3
4ebc27c3
00070aa7
7c0c4c74
4c946007
001c40d7
26e4ff66
75224834
00a0331c
323c4094
60f70010
14c305c3
36c328c3
0aa1f2bc
35740007
14c305c3
36c328c3
0aa222bc
2d740007
05c3c037
2f3c14c3
60a60080
0ab5cabc
23740007
6ea76097
40d72094
60877522
323c1c94
4f3c0010
343c0140
05c3fc7e
2f3c14c3
36c30100
0aa1f2bc
0d740007
00079f5c
0027af5c
14c305c3
36c327c3
0ac37cbc
04150007
ff74001c
00060053
e0760596
08040f56
3f36f016
d0c39696
4177b1c3
7d97c3c3
0f546027
07d46027
901c63c3
60070010
16531154
0b546047
e4dc6067
0193000a
901c63c3
801c0010
01730000
901cc026
86c30020
c02600d3
0010901c
0002801c
10f8a01c
0000a11c
640c1ac3
08068c0c
44c62006
51d4301c
0016311c
70c34664
0007b066
001102dc
32c35e57
0e9460c7
0007cf5c
20773d57
00479f5c
1dc3c0f7
61572bc3
0b09e6bc
5e570233
60a732c3
cf5c0f94
3d570007
9f5c2077
c0f70047
2bc31dc3
10bc6157
50c30b07
5e570d13
618732c3
3b3c5794
61120010
01804f3c
331c2006
15f40100
640c1ac3
20068c4c
301c44c6
311c51d4
46640016
ff51501c
40061a53
3dc3500d
702d6ca2
80452025
080c213c
f6741be4
1a801f3c
20066500
f385135c
1f3c4025
65001a80
135c2006
423cf385
af3c0010
cf5c0180
5d570007
9f5c4077
c0f70047
61376026
1ac307c3
615724c3
0b09d2bc
831c50c3
1f540002
0007cf5c
40775d57
60b76106
2046c0f7
1e972137
24c31ac3
d2bc6157
b4000b09
2ac301d3
8c4c680c
44c62006
51d4301c
0016311c
501c4664
10b3ff7b
4e94a007
0001831c
831c2854
57540002
400728c3
7e576294
20c713c3
273c0654
13c30080
02942187
601c5e97
611c10fc
780c0000
01808f3c
08c38dcc
602617c3
50c34664
2c940007
8e0c780c
3dd708c3
7e1721c3
09534664
32c35e57
075460c7
0180273c
31c33e57
02946187
601c5e97
611c10fc
780c0000
01808f3c
08c38e4c
602617c3
50c34664
780c0bf2
08c38e8c
21c33dd7
46647e17
000750c3
301c2754
311c10f8
6c0c0000
07c38c4c
44c62006
51d4301c
0016311c
04f34664
01804f3c
17c304c3
44bc29c3
04c30aa1
21c33dd7
9ebc7e17
01530aa1
10f8301c
0000311c
8c4c6c0c
15c307c3
301cf073
311c10f8
6c0c0000
07c38c4c
44c62006
51d4301c
0016311c
a0064664
6a9605c3
0f56fc76
00000804
3f36f016
50c3f396
c2c371c3
2006d3c3
21b72337
03004f3c
02806f3c
26c314c3
22bc37c3
00070aa2
001563dc
02c08f3c
05c3e037
28c314c3
88bc6026
00070ab8
0014a3dc
75004317
fff1035c
fff9135c
01c02f3c
02403f3c
0aa2d6bc
ff66201c
b3dc0007
62570013
199460c7
14c305c3
37c326c3
0aa222bc
d3dc0007
e0370012
14c305c3
616628c3
0ab888bc
33dc0007
62d70012
0294331c
0011e4dc
0300af3c
1ac305c3
02802f3c
22bc37c3
00070aa2
001123dc
b53c6317
b31c309d
b4dc0004
60250010
05c36337
2f3c1ac3
37c30200
0aa1f2bc
f3dc0007
6217000f
b6dc6807
901c000f
911c10f8
29c30000
8c0c680c
20060806
301c44c6
311c51c0
46640016
506660c3
92dc0007
6317000e
42173580
08cbb0bc
22176317
63376c80
1ac305c3
01802f3c
0aa282bc
06150007
640c19c3
06c38c4c
29c30f13
8c0c680c
20060806
301c44c6
311c51c0
46640016
0ef280c3
640c19c3
06c38c4c
44c618c3
51c0301c
0016311c
50664664
62571713
3a9460c7
05c3e037
2f3c1ac3
3bc302c0
0ab888bc
0f150007
680c29c3
06c38c4c
44c62006
51c0301c
0016311c
19c34664
0833640c
1f3c02d7
08bc01c0
00070aa3
63172b74
602555a2
40876337
05c32594
03001f3c
02802f3c
f2bc37c3
00070aa1
08c31b74
35004317
b0bc4297
631708cb
6c802297
63176337
602555a2
40876337
05c30b94
03001f3c
02802f3c
f2bc37c3
00070aa1
501c1a15
511c10f8
740c0000
06c38c4c
44c62006
51c0301c
0016311c
740c4664
08c38c4c
44c62006
51c0301c
0016311c
0a334664
40374197
607761d7
74802317
429760b7
625740f7
8f5c6137
0cc300a7
26c31dc3
a6bc6217
701c0ac4
711c10f8
00070000
7c0c1815
06c38c4c
44c62006
51c0301c
0016311c
7c0c4664
08c38c4c
44c62006
51c0301c
0016311c
201c4664
0473ff66
8c4c7c0c
200606c3
301c44c6
311c51c0
46640016
8c4c7c0c
200608c3
301c44c6
311c51c0
46640016
431705c3
42973500
08cbb0bc
229705c3
0ab8c4bc
007320c3
ff74201c
0d9602c3
0f56fc76
00000804
3f36f016
80c3f996
a2c341c3
213c61b7
313c0010
663203f0
333c69a0
62320037
15c3a006
ff53001c
c80c4197
37e476c3
000809dc
08c31173
d184d8c3
4c093dc3
0010313c
602521a2
b33c01a2
78c30010
dda23bc3
74544007
76354547
74352547
72350547
7035c547
6eb44f47
6cb42f47
6ab40f47
68b4cf47
fd50323c
69a22cc3
313c6077
69a2fd50
400660b7
055407a7
fd50303c
5da27cc3
c7a7e006
763c0554
1cc3fd50
6097e7a2
20576432
11ac313c
1f5c6177
3ac300a1
a0252ea1
0c5407a7
108c323c
103c0097
213721ac
00813f5c
66a11ac3
c7a7a025
1b3c3354
323c0010
60f733ac
00617f5c
faa16ac3
80079f85
08c31e54
640760a2
61a70554
61470354
20251694
2dc39fe5
68890093
9fe52025
83d24025
fa546407
079461a7
14548007
68a228c3
9fe52025
0e946147
00b3a025
5258c01c
0016c11c
e5dc8067
0197fff7
0006a00f
001c0073
0796ff66
0f56fc76
00000804
0736f016
52c3ff96
9f5c83c3
12640164
2037cc0c
47f24297
5218301c
0016311c
60376ca2
19940027
00013f5c
65673064
67a70654
61470954
01731094
10c36066
42c34006
606601f3
20c32006
015341c3
20066066
00b321c3
60260006
20c310c3
a3c340c3
6257a684
a7e473c3
301c0635
79c3ff7c
2e54e007
163c0cf2
31c30010
000709c3
2f5c2494
57210001
03f331c3
0030363c
e00779c3
04a61a94
363c1721
27d20010
55a14646
e8466025
01d3f5a1
066647d2
602515a1
55a14886
87d200f3
f5a1e606
08266025
602515a1
680f28c3
03c36006
e0760196
08040f56
3f36f016
02b7f296
82c351c3
9f5c73c3
213c0324
60660020
3230141d
100c133c
03f0313c
308c233c
0001931c
223c0494
01130037
0026393c
0b0d333c
7f5233c4
e0072383
001142dc
83778006
0b0d383c
633c7fe5
2880f88c
5c0c2337
043512e4
52dcc007
af5c0010
b01c0144
dbc30000
3ac30eb3
c35c8c09
2c490009
b21c22f7
343c0003
6277108c
20373c0c
40774006
09c3c0b7
01213f5c
28c313c3
03403f3c
0ac812bc
5d940007
0034343c
208c2c3c
212c133c
5c0c2237
00774037
09c3c0b7
01013f5c
28c313c3
03403f3c
0ac812bc
47940007
00f43c3c
463242d7
112c133c
5c0c21f7
00774037
09c3c0b7
00e13f5c
28c313c3
03403f3c
0ac812bc
31940007
14c382d7
003f141c
5c0c21b7
00774037
09c3c0b7
00c13f5c
28c313c3
03403f3c
0ac812bc
1d940007
931cbfa5
14540002
0001d21c
00f43d3c
aed26ff2
20373c0c
40774026
09c3c0b7
28c32146
03403f3c
0ac812bc
a21c06f2
a0470003
00068bb4
6254a007
60940007
a04740c3
80260294
2bc32297
209da13c
85d254c3
31c32297
ac293b84
108c3a3c
bf3c6177
3c0c0340
40062037
c0b74077
3f5c09c3
13c300a1
3bc328c3
0ac812bc
3e940007
208c353c
00342a3c
21aca23c
0087af5c
20373c0c
c0b70077
2f5c09c3
12c30081
3bc328c3
0ac812bc
28940007
8fd25c0c
00f4353c
100ca33c
0067af5c
00774037
09c3c0b7
00612f5c
00f312c3
60264037
c0b76077
27a609c3
3bc328c3
0ac812bc
9c0c0df2
20268037
c0b72077
27a609c3
3f3c28c3
12bc0340
00070ac8
931c1094
0d540002
60377c0c
80778026
09c3c0b7
28c32146
03403f3c
0ac812bc
23176357
32e421c3
931c0854
05540001
001c04f2
0133ff66
07f27c0f
001cc6d2
0073ff36
ff53001c
fc760e96
08040f56
ff961016
80378006
0ac880bc
08560196
00000804
ff961016
80378026
0ac880bc
08560196
00000804
ff961016
80378046
0ac880bc
08560196
00000804
0336f016
62c3fb96
000753c3
40075a54
60075854
20275654
6c0c1b94
18546007
03c36009
00f71a05
00610f5c
4cb406c7
51e0301c
0016311c
61376c22
00ff331c
2f5c4354
580d0081
0006340f
413c07f3
80070014
213c3694
740c088c
311432e4
701c24c3
711c51e0
04d30016
43c36009
80b79a05
00414f5c
0009905c
24b486c7
fd00893c
00278f5c
00213f5c
1cb466c7
973c9e22
0045309d
00ff431c
931c1554
125400ff
24ac843c
00078f5c
00013f5c
40257921
20073fc5
540fda94
00d301c3
ff53001c
001c0073
0596ff66
0f56c076
00000804
0736f016
80c3fe96
42c361c3
000753c3
40073f54
60073d54
313c3b54
733c080c
740c0010
400612c3
2a3437e4
38c30633
a03c0d22
9a3c208c
39c30300
00079f5c
0039931c
93c30635
0007921c
00079f5c
00f4303c
0300933c
9f5c09c3
931c0027
06350039
921c90c3
9f5c0007
0f5c0027
040d0001
00213f5c
4025642d
26e42045
0006d714
669d043c
0006f40f
001c0073
0296ff53
0f56e076
00000804
01c330c3
023513e4
080403c3
606f6006
080460ef
4006f016
31350087
0a9462bc
401c50c3
411c10fc
700c0000
101c6d8c
111caaab
36643eaa
900c70c3
05c3d18c
0a9404bc
366471ac
0bfd1cbc
aaab101c
3f2a111c
40c36664
101c07c3
111c999a
2cbc4019
14c30a95
0a952cbc
111c2006
08bc40a0
7ebc0a95
20c30a7c
0f5602c3
00000804
0136f016
41c350c3
73c362c3
00c48f5c
3b540007
39542007
37546007
35544007
600738c3
64093254
dfe563f2
7c098025
821c64f2
e025ffff
5ebc05c3
52460ae2
25940007
14c305c3
e8bc26c3
00070ae4
453c1694
04c30100
0ae25ebc
05c306d2
0ae27ebc
02735246
17c304c3
e8bc28c3
20c30ae4
04c30cd2
0ae27ebc
7ebc05c3
201c0ae2
0073ff62
ff53201c
807602c3
08040f56
40c31016
0ae27ebc
0100043c
0ae27ebc
08040856
0f36f016
90c3f296
b2c3a1c3
6f3c83c3
5f3c0280
7f3c0180
60060080
60776037
15c306c3
a4bc27c3
92460ae2
34940007
18c306c3
e8bc45d7
00070ae4
05c31994
46572617
0ae4e8bc
12940007
16c305c3
37c329c3
0afbd4bc
00079206
07c31194
60bc1ac3
50c30af2
0af291e6
92260073
07c300f3
0ae318bc
0c0f3bc3
0f3c45c3
7ebc0080
0f3c0ae2
7ebc0180
0f3c0ae2
7ebc0280
04c30ae2
f0760e96
08040f56
0736f016
70c3f696
92c381c3
5f3ca3c3
6f3c0180
60060080
60776037
16c305c3
a4bc23c3
92460ae2
27940007
18c305c3
e8bc29c3
92260ae4
17940007
0100073c
27c315c3
d4bc36c3
92060afb
06c30ef2
60bc1ac3
50c30af2
07f291e6
18bc06c3
64970ae3
45c30c0f
00800f3c
0ae27ebc
01800f3c
0ae27ebc
0a9604c3
0f56e076
00000804
0136f016
71c3ff96
83c362c3
0ae318bc
a4e640c3
0200031c
031c3154
0eb40200
031ca3a6
2a540100
031ca446
26540180
031ca2a6
16940080
a5c60433
0300031c
031c1d54
06b40300
031ca546
0a940280
a62602b3
0380031c
a6861154
0400031c
043c0d54
9cbc180c
303c0aca
04c3e88b
0010133c
0aca92bc
07c350c3
25c316c3
0b1bf6bc
58090bf2
351c32c3
6037000c
00012f5c
38c3580d
0196ac0f
0f568076
00000804
ff967016
62c350c3
babc43c3
0af20acb
4197700c
05c34037
23c316c3
78bc6157
01960acb
08040e56
01c330c3
023513e4
080403c3
428f5fe6
42af4006
40ef406f
41ef416f
0804426f
50c33016
26bc41c3
96af0acc
0c560006
00000804
3f36f016
c0c3e696
92c361c3
bf3cd3c3
af3c0580
5f3c0480
a0370180
00808f3c
00278f5c
1ac30bc3
03802f3c
02803f3c
0ae2a4bc
00079246
000984dc
16c305c3
e8bc4286
00070ae4
08c32d94
0140163c
e8bc4286
00070ae4
61972594
32dc6007
60970008
7f546007
0100793c
17c305c3
0ae542bc
77941fe7
17c308c3
0ae542bc
71941fe7
1cc30ac3
e8bc4286
0af20ae4
17c308c3
b8bc2bc3
91260afb
47940007
92260073
0ac30893
27c31bc3
74bc3ac3
91660af5
3b940007
0180af3c
03808f3c
1f3c0ac3
27c30580
74bc38c3
00070af5
5f3c2e94
093c0480
15c30200
35c329c3
0afbd4bc
000780a5
093c2294
18c30300
38c329c3
0afbd4bc
19940007
02806f3c
18c305c3
36c329c3
0af574bc
0ff29166
17c306c3
26bc26c3
50c30af5
0ac308f2
42bc16c3
45c30ae5
02d24026
3dc34006
0f3c4c0f
7ebc0080
0f3c0ae2
7ebc0180
0f3c0ae2
7ebc0480
0f3c0ae2
7ebc0380
0f3c0ae2
7ebc0580
0f3c0ae2
7ebc0280
00730ae2
fc7390e6
1a9604c3
0f56fc76
00000804
40c31016
6027628c
08050494
0ae27ebc
0300043c
0ae27ebc
0200043c
0ae27ebc
0100043c
0ae27ebc
7ebc04c3
08560ae2
00000804
3f36f016
0137e296
62c320f7
723c43c3
07c30100
0ae318bc
028630c3
20bc13c3
90c30acc
0140cf3c
1cc304c3
f6bc29c3
40c30b1b
54dc0007
2f5c000b
32c300a1
000c351c
2f5c60b7
2f5c0041
5f3c00a5
df3c0680
8f3c0580
af3c0480
bf3c0380
bf5c0280
00770007
1dc305c3
3ac328c3
0ae2a4bc
00079246
000944dc
1cc305c3
e8bc29c3
92260ae4
77940007
202605c3
0ae55abc
00279106
05c37094
2dc317c3
0afbb8bc
00079126
063c6894
15c30200
38c326c3
0afbd4bc
00079206
08c35e94
28c317c3
0af526bc
00079146
0bc35694
42862117
0ae4e8bc
000780e5
063c4e94
18c30400
aabc2ac3
91860aef
45940007
1bc30ac3
7abc2ac3
80250ae6
3d940007
03805f3c
1f3c05c3
27c30580
74bc35c3
91660af5
31940007
60076497
63972d54
2a546007
04800f3c
0ae318bc
05c340c3
0ae318bc
20d750c3
600600b3
00df313c
82678025
0f3cfbf4
60bc0480
91e60af2
13940007
13c360d7
05c32285
400600b3
00df213c
02670025
0f3cfbf4
60bc0380
40c30af2
90e60053
02800f3c
0ae27ebc
03800f3c
0ae27ebc
04800f3c
0ae27ebc
05800f3c
0ae27ebc
06800f3c
0ae27ebc
1e9604c3
0f56fc76
00000804
60c37016
42c351c3
05d42007
ff53001c
28f44007
24d4a847
0006782c
22547fe7
60d4301c
0016311c
01934006
06f48007
01c32c2c
049440e4
51e40113
402506f4
2c0c6685
019334f2
323c582f
101c0347
111c60d4
6c800016
0006784f
001c0073
0e56ff56
00000804
02d230c3
03c3600c
00000804
400c0bd2
13e432c3
20070715
606c0574
1a1d033c
00060053
00000804
ff961016
60d4301c
0016311c
00534006
133c4025
20371a4f
4f5c3cf2
34c30001
02741fe7
20066026
021502e4
31832026
0014033c
08560196
00000804
50c33016
ff53301c
18bc0dd2
40c30ace
08f26006
0100053c
0ace18bc
02f234c3
03c36026
08040c56
ff53301c
600609d2
602f604f
614f60cf
624f61cf
03c3226f
00000804
5fc62006
0ace5ebc
00000804
03d230c3
6c0c604c
080403c3
0ace72bc
05f40007
0050303c
080c033c
00000804
40c37016
52c361c3
ff53001c
30548007
60d4201c
0016211c
04b32006
4685696c
209434e4
313caad2
201c0347
211c60d4
6d000016
140f0d4c
313ccad2
201c0347
211c60d4
6d000016
180f0d2c
00d7313c
0010233c
60d4301c
0016311c
2a1d033c
202500f3
6007680c
001cda94
0e56ff52
00000804
1f36f016
50c3fe96
b2c3a1c3
0007c3c3
20074b54
40074954
60074754
20064554
e4bc4317
40c30acd
40940007
00c0653c
01c0753c
02c0853c
03c0953c
00770037
17c306c3
39c328c3
0ae2a4bc
00079066
06c32d94
42061ac3
0aee3abc
000740c3
07c31694
42061bc3
0aee3abc
0ff240c3
202608c3
0ae56cbc
740f6046
1cc309c3
3abc4206
40c30aee
10540007
7ebc06c3
07c30ae2
0ae27ebc
7ebc08c3
09c30ae2
0ae27ebc
401c0073
04c3ff53
f8760296
08040f56
0f36f016
80c3fe96
a2c391c3
e2d7b3c3
38540007
36542007
34544007
32546007
3054e007
60d4501c
0016511c
0253c006
07c3944c
08920ebc
00770364
17c304c3
00213f5c
2abc23c3
01640892
08d2a685
740cc025
ed946007
ff74001c
363c02b3
233c00d7
301c0010
311c60d4
133c0016
20372a1d
19c308c3
3bc32ac3
0acebcbc
001c0073
0296ff53
0f56f076
00000804
ff961016
803780d7
0acebcbc
08560196
00000804
50c37016
000761c3
7ebc1954
053c0ae2
7ebc0100
053c0ae2
7ebc0200
301c0ae2
311c10f8
6c0c0000
05c38c4c
44a616c3
631c301c
0016311c
0e564664
00000804
68bc2006
08040acf
0736f016
70c3f696
92c381c3
0007a3c3
20073b54
40073954
60073754
5f3c3554
6f3c0180
60060080
60776037
16c305c3
a4bc23c3
40c30ae2
28940007
17c305c3
3abc4206
40c30aee
15940007
18c306c3
3abc4206
40c30aee
09c30ef2
25c31ac3
d2bc36c3
40c30ab9
619706f2
609763d2
90e662f2
01800f3c
0ae27ebc
00800f3c
0ae27ebc
401c0073
04c3ff56
e0760a96
08040f56
1f36f016
70c3fd96
52c361c3
02d2c3c3
401c44f2
0c13ff53
0014313c
ff56401c
5a546007
00c0823c
01c0923c
02c0a23c
03c0b23c
20372006
08c32077
2ac319c3
a4bc3bc3
40c30ae2
906603d2
7c0908b3
07546087
05546047
03546067
ff74401c
ffe0233c
3f5c40b7
60270041
80072735
363c2794
633cfff0
05c3088c
2cc316c3
0acde4bc
402640c3
0007540f
08c31994
26c33d00
0ae4e8bc
000740c3
363c1194
09c30010
26c33d80
0ae4e8bc
08f240c3
20260ac3
0ae56cbc
401c01f3
08c3ff52
0ae27ebc
7ebc09c3
0ac30ae2
0ae27ebc
7ebc0bc3
04c30ae2
f8760396
08040f56
d6bc6006
08040acf
50c37016
811761c3
13c302c3
46bc24c3
0af20ad0
404634c3
1e7f233c
15c303c3
e8bc26c3
0e560ae4
00000804
0336f016
70c3fd96
02c351c3
e00763c3
60074b54
40074954
2cbc4774
00070ace
353c4354
60070014
863c3f54
963c0100
40060200
40774037
18c306c3
600629c3
0ae2a4bc
03d240c3
07939066
60877c09
60470754
60670554
401c0354
133cff74
20b7ffe0
00413f5c
21356027
21948007
fff0353c
088c533c
173c06c3
25c30010
0ae4e8bc
000740c3
353c1494
08c30010
25c33d80
0ae4e8bc
0bf240c3
202609c3
0ae56cbc
401c01f3
0193ff56
ff52401c
7ebc06c3
08c30ae2
0ae27ebc
7ebc09c3
04c30ae2
c0760396
08040f56
fe96f016
701c60c3
711c10f8
7c0c0000
06068c0c
44a616c3
6330301c
0016311c
50c34664
1e540007
46062006
0891b0bc
746f6006
756f74ef
60776037
153c05c3
253c0100
a4bc0200
0cd20ae2
8c4c7c0c
16c305c3
301c44a6
311c6330
46640016
05c3a006
0f560296
00000804
c6bc0006
08040ad0
60c3f016
42c371c3
27540007
25542007
23544007
2cbc002c
301c0ace
0007ff56
784c1e54
700cac0c
053435e4
301cb00f
02b3ff7c
07c3b00f
25c32006
0891b0bc
03c0463c
18bc04c3
74200ae3
3d8004c3
0af260bc
007330c3
ff53301c
0f5603c3
00000804
40c33016
02d251c3
001c24f2
0233ff53
0ae542bc
043c0ef2
153c0100
42bc0100
07f20ae5
0200043c
0200153c
0ae542bc
08040c56
0f36f016
70c3ff96
92c3a1c3
0b0d313c
233c7fe5
4037f88c
4cd20dd2
6ad239c3
6c0c604c
60256112
640f19c3
ff36501c
e0070fb3
40177954
76944007
600739c3
1c2c7354
0ace2cbc
6e540007
0c107c4c
080c383c
0010b33c
640c19c3
05343be4
501c6411
0c53ff7c
3ac32086
301c2c0d
311c10f8
6c0c0000
001c8c0c
20170100
301c44c6
311c62dc
46640016
b06660c3
4c540007
00012f5c
201c12c3
b0bc0100
473c0891
04c300c0
0ae318bc
642018c3
398004c3
0af260bc
000750c3
0a3c2694
16c30010
b0bc28c3
06c308cb
00012f5c
201c12c3
b0bc0100
473c0891
04c301c0
0ae318bc
642018c3
398004c3
0af260bc
0bf250c3
0010383c
09802ac3
28c316c3
08cbb0bc
6c1139c3
10f8301c
0000311c
8c4c6c0c
200606c3
301c44c6
311c62dc
46640016
501c0073
05c3ff56
f0760196
08040f56
401c1016
64f2ff52
0ad14cbc
04c340c3
08040856
0f36f016
40c3ff96
b2c381c3
000793c3
0009c3dc
0ace2cbc
72dc0007
3b3c0009
7fe50b0d
f88c133c
28c32037
15544007
13542007
600739c3
343c1054
101c0347
111c60d4
6c800016
61126c0c
29c36025
501c680f
0f73ff36
600738c3
20177654
73942007
400729c3
343c7054
101c0347
111c60d4
6c800016
373cec0c
a33c080c
680c0010
06343ae4
4c1139c3
ff7c501c
40860bd3
440d1bc3
10f8301c
0000311c
8c0c6c0c
0100001c
44c62017
62f0301c
0016311c
60c34664
0007b066
3f5c4854
13c30001
0100201c
0891b0bc
18bc08c3
7c200ae3
398008c3
0af260bc
000750c3
0b3c2594
16c30010
b0bc27c3
06c308cb
00012f5c
201c12c3
b0bc0100
483c0891
04c30100
0ae318bc
04c37c20
60bc3980
50c30af2
373c0bf2
1bc30010
16c30580
b0bc27c3
29c308cb
301c4811
311c10f8
6c0c0000
06c38c4c
44c62006
62f0301c
0016311c
00734664
ff56501c
019605c3
0f56f076
00000804
40c33016
02d251c3
001c24f2
0233ff56
0ae35abc
043c0ef2
153c0100
5abc0100
07f20ae3
0200043c
0200153c
0ae35abc
08040c56
40c31016
10540007
7ebc0185
043c0ae2
7ebc01c0
043c0ae2
7ebc02c0
043c0ae2
36bc03c0
08560afd
00000804
0736f016
50c3f596
a2c361c3
24f202d2
ff56401c
301c1233
311c10f8
6c0c0000
36646d2c
3f5c00b7
43c30041
42dc6007
953c0008
09c30200
5abc2006
40c30ae5
05c30ff2
6cbc14c3
053c0ae5
14c30100
0ae56cbc
202609c3
0ae56cbc
8f3c0db3
7f3c01c0
600600c0
60776037
17c308c3
a4bc23c3
90660ae2
5e940007
16c309c3
4ebc2ac3
40c30ae8
4e940007
16c309c3
b8bc28c3
40c30afb
46940007
17c308c3
0af0f6bc
000740c3
07c33f94
27c316c3
0af526bc
000740c3
08c33794
28c317c3
0aefaabc
000740c3
7f3c2f94
07c301c0
27c316c3
0af526bc
000740c3
05c32594
00c01f3c
aabc25c3
40c30aef
1c940007
16c305c3
4ebc2ac3
40c30ae8
14940007
05c3a205
25c317c3
0aefaabc
0cf240c3
16c305c3
4ebc2ac3
40c30ae8
09c305f2
6cbc2026
0f3c0ae5
7ebc01c0
0f3c0ae2
7ebc00c0
04c30ae2
e0760b96
08040f56
0f36f016
70c3f696
83c391c3
0264bf5c
92dc0007
2007001b
001b62dc
32dc6007
af3c001b
40060180
40774037
1f3c0ac3
32c30080
0ae2a4bc
000740c3
001a64dc
0100693c
19c307c3
0ae35abc
000740c3
073c4694
16c30100
0ae35abc
000740c3
593c3e94
073c0200
15c30200
0ae35abc
000740c3
05c33494
f6bc1ac3
40c30af0
2d940007
18c30ac3
4ebc2bc3
40c30ae8
25940007
16c305c3
aabc25c3
40c30aef
1d940007
18c305c3
4ebc2bc3
40c30ae8
15940007
15c305c3
7abc25c3
40c30ae6
68940007
18c305c3
0ae542bc
09541fe7
18c305c3
98bc25c3
40c30ae6
5a948007
00805f3c
1f3c09c3
25c30180
0ae698bc
000740c3
05c34f94
5abc14c3
1fe70ae5
05c30994
25c318c3
0ae67abc
000740c3
5f3c4194
05c30180
25c319c3
0ae67abc
000740c3
05c33794
42bc18c3
1fe70ae5
05c30954
25c318c3
0ae698bc
000740c3
7f3c2994
5f3c0180
07c30080
25c315c3
0aefaabc
000740c3
05c31d94
2bc318c3
0ae84ebc
000740c3
05c31594
27c315c3
0ae67abc
000740c3
07c36c94
42bc18c3
1fe70ae5
07c30954
27c318c3
0ae698bc
800740c3
5f3c5e94
05c30180
00801f3c
7abc25c3
40c30ae6
53940007
18c305c3
0ae542bc
09541fe7
18c305c3
98bc25c3
40c30ae6
45940007
16c306c3
7abc26c3
40c30ae6
3d940007
18c306c3
0ae542bc
09541fe7
18c306c3
98bc26c3
40c30ae6
2f940007
16c306c3
0af0f6bc
000740c3
06c32894
2bc318c3
0ae84ebc
000740c3
5f3c2094
06c30080
f6bc15c3
40c30af0
17940007
18c305c3
4ebc2bc3
40c30ae8
4d940007
60076097
61570ef4
341c6c0c
69d20001
18c305c3
7abc25c3
40c30ae6
3d948007
00800f3c
94bc10c3
40c30ae5
35940007
19c306c3
aabc26c3
40c30aef
2d940007
18c306c3
4ebc2bc3
40c30ae8
25940007
01800f3c
f6bc19c3
40c30af0
1d940007
18c309c3
4ebc2bc3
40c30ae8
15940007
16c309c3
98bc29c3
40c30ae6
60940007
14c309c3
0ae55abc
09941fe7
18c309c3
7abc29c3
40c30ae6
52948007
16c309c3
98bc29c3
40c30ae6
4a940007
14c309c3
0ae55abc
09941fe7
18c309c3
7abc29c3
40c30ae6
3c940007
19c306c3
98bc26c3
40c30ae6
34940007
14c306c3
0ae55abc
09941fe7
18c306c3
7abc26c3
40c30ae6
26940007
1f3c06c3
26c30180
0aefaabc
000740c3
06c31d94
2bc318c3
0ae84ebc
000740c3
06c31594
00801f3c
98bc26c3
40c30ae6
06c30df2
5abc14c3
1fe70ae5
06c30794
26c318c3
0ae67abc
0f3c40c3
7ebc0180
0f3c0ae2
7ebc0080
00730ae2
ff56401c
0a9604c3
0f56f076
00000804
3f36f016
50c3f596
62c3b1c3
9f5c83c3
cf5c02c4
000702e4
002b32dc
02dc2007
4007002b
002ad2dc
400729c3
002a92dc
0394b6e4
56c3b0c3
10f8301c
0000311c
8ccc6c0c
1bc305c3
39c326c3
00b74664
00413f5c
600743c3
002a32dc
01c07f3c
40374006
07c34077
00c01f3c
a4bc32c3
40c30ae2
44dc0007
db3c0029
09c30100
27c31dc3
0ae698bc
000740c3
002704dc
1bc305c3
0ae542bc
54dc0007
4b3c0027
04c30200
0ace18bc
d2dc0007
053c0026
14c30200
0ae542bc
54dc0007
453c0026
04c30100
42bc1dc3
08d20ae5
17c304c3
0ae542bc
74dc0007
0f3c0025
7ebc01c0
0f3c0ae2
7ebc00c0
cf5c0ae2
05c30007
28c316c3
6cbc39c3
40c30ad3
053c4a33
18c30100
0ae35abc
000740c3
053c5494
1ac30200
0ae35abc
000740c3
000a64dc
02005b3c
18bc05c3
00070ace
7f3c4654
05c301c0
f6bc17c3
40c30af0
54dc0007
07c30009
2cc319c3
0ae84ebc
000740c3
0008c4dc
16c307c3
aabc26c3
40c30aef
34dc0007
06c30008
2cc319c3
0ae84ebc
000740c3
05c37a94
27c317c3
0aefaabc
000740c3
07c37294
2cc319c3
0ae84ebc
000740c3
0f3c6a94
18c301c0
aabc28c3
40c30aef
61940007
19c308c3
4ebc2cc3
40c30ae8
59948007
01c05f3c
15c30ac3
0af0f6bc
000740c3
05c35094
2cc319c3
0ae84ebc
000740c3
7f3c4894
0bc300c0
27c315c3
0aefaabc
000740c3
07c33e94
2cc319c3
0ae84ebc
000740c3
0ac33694
25c315c3
0aefaabc
000740c3
05c32e94
2cc319c3
0ae84ebc
000740c3
0dc32694
25c315c3
0aefaabc
000740c3
05c31e94
2cc319c3
0ae84ebc
000740c3
08c31694
28c315c3
0ae698bc
000740c3
001214dc
14c308c3
0ae55abc
0a941fe7
19c308c3
7abc28c3
40c30ae6
24dc8007
5f3c0011
05c301c0
25c315c3
0ae67abc
000740c3
001074dc
19c305c3
0ae542bc
0a541fe7
19c305c3
98bc25c3
40c30ae6
84dc0007
5f3c000f
05c301c0
25c318c3
0ae67abc
000740c3
000ed4dc
19c305c3
0ae542bc
0a541fe7
19c305c3
98bc25c3
40c30ae6
e4dc0007
06c3000d
00c01f3c
98bc26c3
40c30ae6
44dc0007
06c3000d
5abc14c3
1fe70ae5
06c30a94
26c319c3
0ae67abc
000740c3
000c54dc
00c05f3c
15c305c3
7abc25c3
40c30ae6
a4dc0007
05c3000b
42bc19c3
1fe70ae5
05c30a54
25c319c3
0ae698bc
000740c3
000ab4dc
00c05f3c
16c305c3
7abc25c3
40c30ae6
04dc0007
05c3000a
42bc19c3
1fe70ae5
05c30a54
25c319c3
0ae698bc
000740c3
000914dc
02004b3c
18bc04c3
00070ace
0ac31254
2ac314c3
0aefaabc
000740c3
000814dc
19c30ac3
4ebc2cc3
40c30ae8
78940007
16c30ac3
aabc2ac3
40c30aef
70940007
19c30ac3
4ebc2cc3
40c30ae8
68940007
01c07f3c
16c307c3
aabc27c3
40c30aef
5e940007
19c307c3
4ebc2cc3
40c30ae8
56940007
16c306c3
0af0f6bc
000740c3
06c34f94
2cc319c3
0ae84ebc
000740c3
5f3c4794
05c300c0
25c316c3
0aefaabc
000740c3
05c33d94
2cc319c3
0ae84ebc
000740c3
07c33594
27c316c3
0aefaabc
000740c3
07c32d94
2cc319c3
0ae84ebc
000740c3
08c32594
f6bc16c3
40c30af0
1e940007
19c306c3
4ebc2cc3
40c30ae8
16940007
1f3c06c3
26c300c0
0ae698bc
000740c3
06c36694
5abc14c3
1fe70ae5
06c30994
26c319c3
0ae67abc
800740c3
5f3c5894
05c300c0
25c316c3
0ae698bc
000740c3
05c34e94
5abc14c3
1fe70ae5
05c30994
25c319c3
0ae67abc
000740c3
5f3c4094
05c300c0
25c316c3
0ae698bc
000740c3
05c33694
5abc14c3
1fe70ae5
05c30994
25c319c3
0ae67abc
000740c3
5f3c2894
05c300c0
25c318c3
0aefaabc
000740c3
05c31e94
2cc319c3
0ae84ebc
000740c3
05c31694
01c01f3c
98bc28c3
40c30ae6
23940007
14c308c3
0ae55abc
09941fe7
19c308c3
7abc28c3
40c30ae6
15948007
6007788c
78ec0df4
341c6c0c
68d20001
19c308c3
7abc28c3
40c30ae6
08c306f2
94bc18c3
40c30ae5
01c00f3c
0ae27ebc
00c00f3c
0ae27ebc
401c0233
01d3ff56
0100863c
0200a63c
16c305c3
0ae35abc
000740c3
ffe0e4dc
04c3b633
fc760b96
08040f56
3f36f016
00f7eb96
92c371c3
df5c60b7
00070404
001d22dc
f2dc2007
4007001c
001cc2dc
20071dc3
001c82dc
02008f3c
200608c3
b0bc4406
301c0891
311c10f8
6c0c0000
40374857
00d78d0c
29c317c3
46643dc3
3f5c0137
43c30081
f2dc6007
0dc3001a
05001f3c
0ae724bc
000740c3
001a64dc
04006f3c
5ebc06c3
40c30ae2
d4dc0007
06c30019
eabc1dc3
40c30aeb
05d250c3
7ebc06c3
32330ae2
c6bc0897
38c30ad0
5b9d033c
13940007
6f3c40c3
00f30200
4a1d063c
68bc2897
80250acf
f97445e4
04000f3c
0ae27ebc
2ef39066
a107a025
0897e494
0ad0c6bc
9066a0c3
3c540007
04005f3c
202605c3
0ae55abc
18940007
1ac307c3
0ae35abc
000740c3
073c2d94
1a3c0100
5abc0100
40c30ae3
24940007
0200073c
02001a3c
0ae35abc
07c30393
2dc315c3
74bc3ac3
40c30af5
14940007
0100073c
2dc315c3
01003a3c
0af574bc
0af240c3
0200073c
2dc315c3
02003a3c
0af574bc
0f3c40c3
7ebc0400
80070ae2
001114dc
60376517
22170ac3
3dc34097
0ad36cbc
000740c3
001054dc
20372517
10c30217
3dc34097
0ad36cbc
000740c3
000f94dc
40374517
10c30217
3dc34097
0ad36cbc
000740c3
000ed4dc
02005f3c
03c06f3c
542c740c
0007df5c
20772517
1ac303c3
36bc6097
40c30ad5
a4dc0007
a085000d
ef9456e4
18bc00d7
103c0ace
21f7fff0
0100393c
293c6177
41b70200
c01c74c3
84c30001
bcc364c3
005354c3
b21ce112
3bc3ffff
21d76ff2
5fe721c3
00d77554
0ace1ebc
61d770c3
3fe513c3
b01c21f7
273c001c
32c30ecb
63f235a3
fcf353c3
0e94a027
25174df2
09c32037
409719c3
6cbc3dc3
40c30ad3
d9540007
c0251333
67202086
300d323c
a04683a3
cf9461e4
c31cc006
21940001
ff80383c
1f3c6212
a5800540
e64e053c
5abc19c3
40c30ae3
7e940007
033c740c
21570100
0ae35abc
000740c3
740c7594
0200033c
5abc2197
40c30ae3
0453c6c3
40374517
19c309c3
3dc34097
0ad36cbc
000740c3
c0256194
f394c087
ff80383c
1f3c6212
65800540
fe64335c
0007df5c
40774517
13c309c3
609729c3
0ad536bc
800740c3
84c34994
a02664c3
0bc3f093
4194a047
3ff4c007
0100ba3c
02007a3c
2cc350c3
65174bf2
09c36037
409719c3
6cbc3dc3
00070ad3
883c2e94
383c080c
60070104
c31c2554
17940001
19c30ac3
0ae35abc
000740c3
0bc31f94
5abc2157
40c30ae3
18940007
219707c3
0ae35abc
11940007
0193c0c3
0007df5c
40774517
1ac309c3
609729c3
0ad536bc
a02504f2
c87456e4
89f240c3
27d22857
1dc309c3
ccbc4517
40c30ad2
28970ac3
0acf68bc
02005f3c
04006f3c
024f053c
68bc2897
56e40acf
0073fa94
ff56401c
159604c3
0f56fc76
00000804
0336f016
60c3fd96
72c391c3
401c83c3
0007ff53
026c2054
0ad0c6bc
906650c3
15540007
6026e037
7a6c6077
08c360b7
00c0163c
39c325c3
0ad80abc
07f240c3
4abc05c3
03f20ace
ff29401c
3a6c05c3
0acf68bc
039604c3
0f56c076
00000804
0336f016
60c3fd96
82c391c3
ff53401c
57540007
c6bc026c
70c30ad0
00079066
784c5054
42062cec
0aee3abc
000740c3
784c4694
0100073c
42062d0c
0aee3abc
000740c3
073c3c94
20260200
0ae56cbc
c6bc1a6c
50c30ad0
00079066
8f5c2754
60260007
7a6c6077
063c60b7
17c303c0
39c325c3
0ad80abc
000740c3
05c31794
00c0163c
0ae542bc
053c0ff2
163c0100
42bc01c0
08f20ae5
0200053c
02c0163c
0ae542bc
401c03d2
05c3ff28
68bc3a6c
07c30acf
68bc3a6c
00730acf
fed3a006
039604c3
0f56c076
00000804
0f36f016
70c3f196
23c362c3
04f2c2d2
ff53501c
06c31e13
0acde4bc
000750c3
000ea4dc
10f8301c
0000311c
8c0c6c0c
15c30946
301c44c6
311c6308
46640016
b06680c3
72dc0007
784c000d
b33c6c0c
07c30080
2bc318c3
0b1bf6bc
000750c3
000b64dc
03c0963c
02c04f3c
00c0af3c
00770037
14c309c3
3f3c2ac3
a4bc01c0
50c30ae2
34dc0007
0037000a
063c0077
163c00c0
263c01c0
35c302c0
0ae2a4bc
000750c3
000944dc
c6bc1a6c
70c30ad0
c2dc0007
784c0008
2c6c04c3
3abc4206
50c30aee
44dc0007
784c0008
2ccc0ac3
3abc4206
50c30aee
7a940007
0f3c784c
2c8c01c0
3abc4206
50c30aee
70940007
07c3784c
42062cec
0aee3abc
000750c3
784c6994
0100073c
42062d0c
0aee3abc
000750c3
073c5f94
20260200
0ae56cbc
18c309c3
e8bc2bc3
50c30ae4
52940007
b0e679ec
4e546007
03c0463c
00c05f3c
15c304c3
0ae542bc
09541fe7
15c304c3
26bc24c3
50c30af5
3c940007
02c03f3c
60266037
5a6c6077
04c340b7
263c17c3
3f3c00c0
0abc01c0
50c30ad8
2a940007
780f6046
3a6c07c3
0acf68bc
01c00f3c
0ae27ebc
02c00f3c
0ae27ebc
00c00f3c
0ae27ebc
284608c3
0b06b8bc
10f8301c
0000311c
8c4c6c0c
200608c3
301c44c6
311c6308
46640016
b06602d3
a007e006
063cb454
7ebc00c0
063c0ae2
7ebc01c0
063c0ae2
7ebc02c0
063c0ae2
36bc03c0
f9330afd
0f9605c3
0f56f076
00000804
3f36f016
a0c3e296
c2c361c3
bf5c93c3
8f5c0524
00070544
000c02dc
40072bc3
000bc2dc
600738c3
000b82dc
400729c3
000b42dc
60073cc3
000b02dc
6047680c
000ac4dc
0c2c39c3
0ace2cbc
54dc0027
5f3c000a
60060580
60776037
1f3c05c3
23c30680
0ae2a4bc
000740c3
000aa4dc
684c29c3
2ccc05c3
3abc4206
40c30aee
24dc0007
05c30008
0ae306bc
363c50c3
30e4180c
303c0535
633c0070
7f3c188c
07c30680
26c31ac3
0ae4e8bc
000740c3
363c6b94
35e4180c
253c7335
07c30074
2d206106
0ae3d4bc
c0250d73
0494c827
ff39401c
29c30ab3
0cc3684c
2f3c2c0c
6c2c0080
0ada84bc
000740c3
0dc34994
2bc315c3
0af526bc
000740c3
2bc34194
6007680c
0dc31094
0ae27ebc
02400f3c
0ae27ebc
03400f3c
0ae27ebc
7ebc07c3
fa930ae2
15c307c3
b8bc27c3
40c30afb
26940007
1bc30ac3
38c325c3
0af574bc
000740c3
0f3c1d94
18c30680
7abc28c3
40c30ae6
14940007
15c308c3
26bc28c3
40c30af5
08c30df2
25c317c3
74bc38c3
40c30af5
28c305f2
6007680c
0f3ca754
b6bc0080
0f3c0ad2
7ebc0580
0f3c0ae2
7ebc0680
02b30ae2
ff56401c
5f3c0253
05c30080
0ace6cbc
ee940007
03c0a93c
df3c60c3
5f3c0140
7f3c0580
f0d30440
1e9604c3
0f56fc76
00000804
1f36f016
70c3f696
82c3a1c3
bf5c93c3
cf5c0284
000702a4
40073454
60073254
3cc33054
2d546007
60073bc3
5f3c2a54
6f3c0180
60060080
60776037
16c305c3
a4bc23c3
40c30ae2
1d940007
c077a037
1ac307c3
3cc32bc3
0adb84bc
08f240c3
19c308c3
36c325c3
0ab9d2bc
0f3c40c3
7ebc0180
0f3c0ae2
7ebc0080
00730ae2
ff56401c
0a9604c3
0f56f876
00000804
84bc6006
08040ada
0736f016
50c3f496
82c371c3
000793c3
0008b2dc
82dc2007
40070008
000852dc
22dc6007
600c0008
14dc6047
002c0008
0ace2cbc
7b540007
2cbc1c2c
00070ace
744c7654
0c4c5c4c
4206284c
08922abc
416440c3
6b948007
c6bc166c
60c30ad0
60f77066
66540007
80778037
02000f3c
01001f3c
34c324c3
0ae2a4bc
000700f7
4f3c4e94
744c0200
2c6c04c3
3abc4206
00f70aee
3b940007
0100af3c
0ac3744c
42062c8c
0aee3abc
000700f7
80373094
40774026
60b7766c
03c0053c
00c0173c
3ac326c3
0ad80abc
000700f7
04c32094
0ae318bc
29c340c3
30e4680c
201c0534
40f7ff7c
08c30293
00613f5c
24c313c3
0891b0bc
18bc06c3
70200ae3
28c306c3
60bc2980
00f70af2
8c0f39c3
01000f3c
0ae27ebc
02000f3c
0ae27ebc
366c06c3
0acf68bc
301c00f3
0073ff53
ff56301c
00d760f7
e0760c96
08040f56
fd961016
80378157
80778197
80b78006
0ad80abc
08560396
00000804
3f36f016
c0c3dd96
d2c3b1c3
af5c93c3
000705e4
001702dc
d2dc2007
40070016
0016a2dc
40074b97
001662dc
60073ac3
001622dc
680f6006
082c2ac3
0ace2cbc
94dc0027
3f3c0015
60370280
03803f3c
0f3c6077
1f3c0780
2f3c0680
3f3c0580
a4bc0480
50c30ae2
00079066
001564dc
00770037
01800f3c
00801f3c
35c325c3
0ae2a4bc
65c304d2
0e1385c3
0e6c3ac3
0ad0c6bc
2ac360c3
c6bc0a6c
80c30ad0
64540007
6254c007
02805f3c
684c2ac3
2ccc05c3
3abc4206
40c30aee
04dc0007
2ac3000f
0f3c684c
2c6c0180
3abc4206
40c30aee
44dc0007
2ac3000e
0f3c684c
2c8c0080
3abc4206
40c30aee
84dc0007
2cc3000d
6007680c
001012dc
680c2bc3
c2dc6007
0cc3000f
42bc15c3
1fe70ae5
000f54dc
15c30bc3
0ae542bc
e4dc1fe7
05c3000e
0ae306bc
393c50c3
30e4180c
303c0535
933c0070
7f3c188c
07c30380
29c31dc3
0ae4e8bc
000740c3
000a94dc
180c393c
49dc35e4
253c000d
07c30074
2d206106
0ae3d4bc
90661973
9f3c1333
0f3c0580
15c30380
39c327c3
0af574bc
000740c3
0008d4dc
0480bf3c
15c30cc3
3bc327c3
0af574bc
000740c3
000814dc
684c2ac3
2cec06c3
3abc4206
40c30aee
76940007
684c2ac3
0100063c
42062d0c
0aee3abc
000740c3
063c6b94
20260200
0ae56cbc
00c00a3c
5abc18c3
40c30ae3
5e940007
01c00a3c
0100183c
0ae35abc
000740c3
0a3c5594
183c02c0
5abc0200
40c30ae3
4c940007
00807f3c
01805f3c
0077a037
16c309c3
37c326c3
0add54bc
000740c3
a0373d94
0bc30077
28c318c3
54bc37c3
40c30add
32940007
01805f3c
1f3c05c3
24bc0880
40c30ae7
28940007
6897a037
08c36077
26c316c3
00803f3c
0ad536bc
000740c3
06c31b94
489715c3
0ad2ccbc
000740c3
5f3c1394
06c30780
02801f3c
26bc25c3
40c30af5
05c309f2
42bc1cc3
04f20ae5
4b976026
06c3680f
2a6c2ac3
0acf68bc
3ac308c3
68bc2e6c
0f3c0acf
7ebc0780
0f3c0ae2
7ebc0680
0f3c0ae2
7ebc0580
0f3c0ae2
7ebc0480
0f3c0ae2
7ebc0280
0f3c0ae2
7ebc0380
0f3c0ae2
7ebc0180
0f3c0ae2
7ebc0080
02730ae2
ff56401c
90e60213
7f3cfa33
5f3c0280
0bc30680
25c317c3
0afbb8bc
000740c3
e593c594
239604c3
0f56fc76
00000804
0736f016
40c3f696
82c391c3
e497a3c3
33540007
31544007
2f54e007
600764d7
60062c54
6f3c7c0f
06c30180
42062006
0891b0bc
00805f3c
200605c3
b0bc4206
04c30891
26c319c3
66bc35c3
40c30abf
e0370bf2
607764d7
15c306c3
3ac328c3
0add62bc
0f3c40c3
7ebc0180
0f3c0ae2
7ebc0080
00730ae2
ff56401c
0a9604c3
0f56e076
00000804
07350047
055400a7
03540087
129400e7
00476406
00471154
620607d4
62860dd2
08940027
68060133
06540087
00a76606
301c0354
03c3ff53
00000804
08040806
01c330c3
023513e4
080403c3
50c33016
1081405c
1a548047
05b48047
802789d2
01b31394
22548087
0e9480a7
103c02f3
48060cc0
0b05a6bc
03f304c3
0cc0103c
2ebc4806
00060b1a
103c0313
48060cc0
0b16f6bc
11540007
103c0273
201c0cc0
f8bc0080
09d20b18
103c0173
201c0cc0
b8bc0080
04f20b19
355c6026
0c56108d
00000804
50c37016
205c61c3
46f21089
0adf5ebc
c4dc0007
355c0009
60471081
60473a54
6bd206b4
e4dc6027
03b30008
6e546087
84dc60a7
09730008
1cc0453c
14c305c3
0b055cbc
153c05c3
480614c0
0b05a6bc
14c305c3
a6bc4206
05c30b05
5cbc16c3
0e130b05
1cc0453c
14c305c3
0b1a6cbc
153c05c3
480614c0
0b1a2ebc
14c305c3
2ebc4286
05c30b1a
6cbc16c3
0b530b1a
1cc0453c
14c305c3
0b173abc
56940007
153c05c3
480614c0
0b16f6bc
4e940007
14c305c3
f6bc4406
00070b16
05c34794
3abc16c3
00070b17
08133d54
1cc0453c
14c305c3
0b187ebc
38940007
153c05c3
201c14c0
f8bc0080
00070b18
05c32f94
460614c3
0b18f8bc
28940007
16c305c3
0b187ebc
1e540007
453c0433
05c31cc0
3ebc14c3
00070b19
05c31994
14c0153c
0080201c
0b19b8bc
10940007
14c305c3
b8bc4806
0af20b19
16c305c3
0b193ebc
600605f2
108d355c
0e560006
00000804
50c3f016
72c361c3
1089305c
5ebc65f2
00070adf
455c2f94
80471081
80471a54
89d205b4
13948027
808701b3
80a71e54
02b30e94
16c305c3
a6bc27c3
04c30b05
05c30333
27c316c3
0b1a2ebc
02530006
16c305c3
f6bc27c3
01930b16
16c305c3
f8bc27c3
00d30b18
16c305c3
b8bc27c3
0f560b19
00000804
2037ff96
205c4006
3f5c108d
305c0001
40171085
604732c3
32c30a35
075460a7
608732c3
32c30454
249460e7
32c34017
17546047
604732c3
4cd205d4
1a944027
401701b3
608732c3
32c31254
129460a7
eebc0173
00170b00
04bc01f3
01930b1a
0b16bebc
1ebc0133
00d30b18
0b17bebc
001c0073
0196ff53
00000804
0336f016
40c3fe96
53c362c3
14c0903c
0ae07ebc
000780c3
000af4dc
10fc301c
0000311c
6c0c6c0c
0bc1035c
035c10c3
203c0bc9
135c40ac
213c0bd1
035c812c
303c0bd9
66d2c12c
ff38001c
59dca1a7
743c0009
345c0cc0
60471081
60472954
6bd205b4
06946027
608702b3
60a74e54
001c3854
1033ff53
1c35a807
16c304c3
a6bc25c3
04c30b05
5cbc17c3
a2060b05
a80701b3
04c30f35
25c316c3
0b1a2ebc
17c304c3
0b1a6cbc
8806a286
a8070973
07c308b4
25c316c3
08cbb0bc
08138806
16c304c3
f6bc25c3
00070b16
04c35694
3abc17c3
a4060b17
00078806
09b33354
0080531c
04c31535
25c316c3
0b18f8bc
43940007
17c304c3
0b187ebc
401ca606
00070080
07331f54
0080531c
07c309b4
25c316c3
08cbb0bc
0080401c
04c30233
25c316c3
0b19b8bc
27940007
17c304c3
0b193ebc
401ca806
04d20080
54e403d3
1e800634
52a02006
0891b0bc
1da26006
161c10c3
2077005c
00210f5c
09a129c3
21c33da2
0036261c
0f5c4037
1da10001
34e46025
08c3ed14
c0760296
08040f56
3f36f016
fddcf21c
a1c300b7
6077b2c3
12849f5c
0adf38bc
601c50c3
0007ff53
000ca3dc
3f5c6026
801c111d
811c10f8
28c30000
8c0c680c
1f5c0806
44c610c4
638c301c
0016311c
70c34664
0007d066
000b22dc
680c28c3
08068c0c
10c41f5c
301c44c6
311c638c
46640016
0ff2c0c3
680c28c3
07c38c4c
10c41f5c
301c44c6
311c638c
46640016
12b3d066
4af24057
07c395c3
00213f5c
25c313c3
0891b0bc
4f3c27c3
04c300c0
39c32097
0ae0bcbc
000760c3
04c36694
2bc31ac3
0ae042bc
000760c3
04c35e94
9abc1cc3
a0c30adf
56940007
9f5cd5c4
8ac31304
0973b4c3
11193f5c
602745c3
80060294
20970bc3
35c32cc3
0ae0bcbc
000760c3
0bc34294
24c317c3
0ae042bc
000760c3
0bc33a94
12a41f5c
12c42f5c
0ae042bc
000760c3
0bc33094
22301f3c
42bc4026
60c30ae0
27940007
17c30bc3
0adf9abc
9d8460c3
1f940007
0e8039c3
58bc15c3
30c30adf
12e42f5c
088402c3
23c317c3
08cbb0bc
3f5c8584
23c31119
40374025
00013f5c
111d3f5c
13042f5c
83e432c3
6ac3b214
10f8501c
0000511c
8c4c740c
1f5c07c3
44c610c4
638c301c
0016311c
740c4664
0cc38c4c
10c41f5c
301c44c6
311c638c
46640016
f21c06c3
fc760224
08040f56
08040046
50c33016
00077fa6
301c1954
311c10f8
6c0c0000
00868c0c
41262006
686c301c
0016311c
146f4664
08d27fc6
600f6006
6026740f
6006742f
03c3744f
08040c56
50c33016
20540007
4006606c
039366f2
103c2006
40252b9d
740c146c
21e413c3
301cf874
311c10f8
6c0c0000
20068c4c
301c4126
311c6860
46640016
746f6006
742f740f
0c56744f
00000804
0736f016
61c350c3
83c372c3
0104af5c
01249f5c
5ebc06d2
40c30ae2
4e940007
06c3c8d2
0ae25ebc
05c340c3
44948007
07c3ebd2
0ae25ebc
06d240c3
7ebc05c3
06c30ae2
38c30733
08c36ed2
0ae25ebc
09d240c3
7ebc05c3
06c30ae2
0ae27ebc
055307c3
60073ac3
0ac31154
0ae25ebc
0cd240c3
7ebc05c3
06c30ae2
0ae27ebc
7ebc07c3
08c30ae2
49c302f3
16548007
5ebc09c3
40c30ae2
10540007
7ebc05c3
06c30ae2
0ae27ebc
7ebc07c3
08c30ae2
0ae27ebc
7ebc0ac3
04c30ae2
0f56e076
00000804
12c3400c
323c4ed2
133c01c7
323cfe40
406c100c
09817f85
20250073
1ef20132
080401c3
0ae306bc
303c4006
62d20074
303c4026
341cf90c
6c000007
09806352
00000804
ff967016
602c50c3
281531e4
0020613c
10f8301c
0000311c
546c6c0c
6848101c
0016111c
8c2c2037
163c02c3
4006100c
46646126
1fc630c3
11546007
542c746f
123cd42f
00d3100c
0006746c
40250ce1
742c2085
20e403c3
0006f874
0e560196
00000804
50c37016
02d241c3
1fa623f2
00060513
255454e4
702c340c
061531e4
28bc04c3
00070ae3
346c1c94
6006506c
613c00d3
623c3a1d
6025027f
60c3140c
f87436e4
000600b3
027f023c
300c6025
36e461c3
140cf974
344c100f
0006304f
08040e56
50c33016
5ebc41c3
05f20ae2
15c304c3
0ae35abc
08040c56
ff961016
3fe531c3
60064180
81a20153
88098037
4f5c81a1
880d0001
3fe56025
31e45fe5
0196f574
08040856
0fd21016
204f2006
406c200f
00b331c3
423c8006
60253b9d
41c3202c
f97434e4
08040856
80261016
313c0093
600ffff0
2007200c
29d203d4
70a00133
333c406c
6981130c
005373d2
0856204f
00000804
51c3f016
323c4026
733c100d
6386fff0
800ccca0
233c6a20
606c130c
40060d00
600c0153
133c2623
21a3508d
fe7f203c
238327c3
80079fe5
0f56f515
00000804
50c37016
200741c3
600c20f4
04d431e4
0ae3acbc
006c0353
100c313c
40062180
313c00d3
303c2a1d
4025027f
6e20740c
f87423e4
600600b3
027f303c
340c4025
fa7421e4
740f6620
08040e56
0136f016
62c351c3
06d42007
acbc06c3
e0060ae3
600c0753
01c7333c
067413e4
5abc16c3
70c30ae3
16c30613
0ae35abc
000770c3
05c32a94
5cbc2386
80c30a7c
05c347c3
6ebc2386
02d20a7c
08c38026
233c7000
00b3100c
85618006
40856025
180c386c
34e440c3
383cf874
2580100c
341d6386
60262530
7fe53223
3083040c
06c3640f
0ae3bebc
807607c3
08040f56
40c37016
200751c3
600c28f4
602c2580
051531e4
0ae328bc
20940007
7500500c
506c700f
621213c3
09807f85
0010353c
333c6ca0
4980130c
00936006
c1e1c981
3fe57f85
fb1515e4
6006106c
203c4006
6025027f
fb7435e4
0e560006
00000804
0136f016
42c351c3
065404e4
5abc14c3
00070ae3
05c34894
5cbc2386
60c30a7c
2180700c
32c3502c
077413e4
202504c3
0ae328bc
37940007
07f4a367
16c304c3
0ae462bc
2f940007
238605c3
0a7c6ebc
000760c3
60262454
833c3023
6386fff0
b06cec20
01c32006
540c0213
600d323c
301c13a3
311cffff
13830fff
027f153c
123c0025
1883708d
02e4500c
27d2ef74
133c706c
323c2b9d
700f0010
bebc04c3
00060ae3
0f568076
00000804
40c37016
52c361c3
6027602c
204606d4
0ae328bc
1c940007
acbc04c3
02530ae3
210604c3
92bc24c3
bfe50ae4
10940007
363c506c
280c009f
680f31a3
6025700c
a007700f
04c3eed4
0ae3bebc
0e560006
00000804
41c31016
045401e4
0ae35abc
600604f2
03c3704f
08040856
800cf016
43e4640c
43e41ad4
343c1a74
233c100c
606cffc0
646ccd00
6006ad00
013323c3
35011901
09b401e4
01e45f85
60250814
f77434e4
00930006
00530026
0f561fe6
00000804
40c37016
a44c604c
36e465c3
361c0a54
333c0001
7fe50b0d
03c37f52
00f30072
03946027
14c301c3
0ae51ebc
08040e56
6027604c
600c0b54
0ad46027
6c0c606c
06b431e4
31e40006
1fe60434
00260053
00000804
50c33016
acbc41c3
746c0ae3
ffff201c
0fff211c
8c0f4283
746c4006
62d26c0c
540f4026
08040c56
20c37016
a38641c3
1150141d
0006600c
091431e4
341d686c
333c2450
32431a1d
0014033c
08040e56
0336f016
41c360c3
702c200c
061531e4
28bc04c3
00070ae3
30102f94
700f780c
621253c3
ffc0233c
83c3786c
706c8284
0006ed00
017310c3
688128c3
088c233c
d92c203c
3f855ce1
0014033c
a007bfe5
500cf415
100c323c
6c80306c
200600b3
027f133c
29e44025
584cfb74
04c3504f
0ae3bebc
c0760006
08040f56
0f36f016
71c350c3
600c62c3
34e4840c
a5c305f4
43c384c3
a1c30073
382c83c3
42e421c3
06c30874
0010143c
0ae328bc
42940007
343c7810
780f0010
3c6c3470
0006b86c
025320c3
2a1d713c
09c36380
2a1d003c
033c6c00
701ce08c
711cffff
37830fff
027f353c
28e44025
84e4ee74
123c1554
0213100c
7c6c7ac3
6380ec81
e08c033c
ffff701c
0fff711c
353c3783
4025027f
24e42085
140ff074
35c3580c
e0060093
4025ec0f
2be46085
06c3fb74
0ae3bebc
f0760006
08040f56
0736f016
71c350c3
041042c3
682cc00c
071536e4
16c304c3
0ae328bc
38940007
d00f3010
5c70b46c
2006106c
025321c3
024f353c
773c7ac3
6fa02a1d
133c6ca0
701cf88c
711cffff
37830fff
027f303c
28e44025
01d3ee74
024f353c
133c6ca0
701cf88c
711cffff
37830fff
027f303c
26e44025
700cf274
e00600b3
027f703c
39e46025
04c3fb74
0ae3bebc
e0760006
08040f56
0136f016
61c370c3
804c52c3
48e40450
884f0594
0ae5d2bc
1ebc01f3
1fe70ae5
14510594
17c306c3
944f0093
16c307c3
30bc25c3
80760ae6
08040f56
0136f016
61c370c3
804c52c3
83c3644c
055448e4
d2bc884f
02730ae5
0ae51ebc
05541fe7
07c3944f
011316c3
0b0d343c
7f327fe5
06c3744f
25c317c3
0ae630bc
0f568076
00000804
50c33016
2007200c
01c31f54
1d542027
1af42027
42c34006
333c746c
001c2a1d
011cffff
30030fff
0b0d333c
7f327fe5
40259180
f17421e4
313c0006
43e4090c
00260474
00060053
08040c56
50c3f016
6007600c
60272054
60272054
06bc1ef4
40c30ae3
20260386
025321c3
62c3746c
1a1d733c
cfd26783
301c4112
311cffff
63c30fff
033526e4
40262025
04e40025
0073ee74
00530006
0f560026
00000804
200c3016
11f42027
4026006c
2a1d303c
ffff401c
0fff411c
35e454c3
40250694
f57421e4
00530026
0c560006
00000804
41c31016
0c0c606c
0014303c
60075fa6
303c1e54
341c0020
61120004
313c2c00
4046028d
133c69a0
313c128d
69a0028d
128d133c
028d313c
333c6d20
201c128d
211cffff
32830fff
4006700f
085602c3
00000804
3f36f016
b0c3fd96
4037a1c3
2077200c
280c2ac3
43c3602c
077414e4
28bc2025
00070ae3
000e94dc
10f8301c
0000311c
8c0c6c0c
1000001c
41262006
682c301c
0016311c
c0c34664
5cc31fc6
42dca007
6bc3000d
2cc3786c
01132006
1a1d033c
8006080f
4105882f
5bc32025
06c3d40c
f57410e4
600600d3
682f680f
20254105
700c4ac3
31e46112
4cc3f715
0000901c
54c308b3
0017700c
23c32006
ffff601c
0fff611c
31c32683
0a7e5abc
00b70683
a8702ac3
0313c006
20060097
233c3dc3
31c36a1d
0a7e5abc
740c81c3
4c00f42c
23e42026
20060214
7c0008c3
540f6580
a105742f
1ac3c025
32c3440c
e57463e4
700c502c
323c7c32
623c21ac
504ce08c
0980b06c
02e42026
20060214
65807700
706f104f
0001921c
5ac38105
06c3d40c
b87490e4
180c393c
c5801cc3
0010593c
180c353c
02f32580
780c582c
323c7c32
823c21ac
440ce08c
8980e42c
42e40026
00060214
7d0028c3
840f6180
2105642f
a025c105
4c0c3ac3
080c323c
53e46025
5bc3e4f4
323c146c
6cc3180c
40063980
313c0173
401c044f
411cffff
34830fff
027f303c
5ac34025
32e4740c
00b3f315
103c2006
4025027f
43c36057
f97424e4
740c5ac3
6bc36025
0bc3780f
0ae3bebc
10f8301c
0000311c
8c4c6c0c
20060cc3
301c4126
311c682c
46640016
1ac30bc3
0ae51ebc
000630c3
06547fe7
1ac30bc3
30bc2bc3
03960ae6
0f56fc76
00000804
3f36f016
81c370c3
a40cc2c3
080c353c
0010433c
01ff431c
531c07d4
04d400ff
0ae74ebc
7c2c0e13
071534e4
14c307c3
0ae328bc
67940007
a01c9c0f
09330000
100c3a3c
8d005c6c
9c3c700c
501c328d
511cffff
95830fff
647018c3
56c3c006
09c30493
3bc32006
6a1d233c
5abc31c3
30c30a7e
300c01c3
20264c80
021423e4
64002006
20260a80
021402e4
45802006
e08c303c
21ac523c
ffff101c
0fff111c
043c0183
c025027f
680c28c3
6de4d3c3
0193d974
7480300c
e08c533c
ffff201c
0fff211c
343c3283
b5f2027f
0001a21c
ac0c38c3
ade4d5c3
07c3b474
0ae3bebc
28c307c3
f4bc280c
07c30ae3
1ebc18c3
30c30ae5
7fe70006
07c30654
27c318c3
0ae630bc
0f56fc76
00000804
4006606c
1000211c
68200c0c
0804640f
3f36f016
70c3ff96
d2c391c3
183c0410
602c080c
051531e4
0ae328bc
4e940007
100cc83c
0010b83c
a4c39c6c
a006ac84
04d365c3
20060dc3
233c3ac3
31c35a1d
0a7e5abc
203730c3
4c00100c
23e42026
20060214
64000017
20260b00
021402e4
65802006
101c20c3
111cffff
21830fff
027f243c
e08c203c
212c633c
58e4a025
d00fda74
34c32bc3
c0060093
4025cc0f
1c0c6085
21e410c3
07c3f974
0ae3bebc
19c307c3
0ae51ebc
07541fe7
19c307c3
30bc27c3
f7330ae6
01960006
0f56fc76
00000804
50c3f016
01c371c3
5cbc2386
40c30a7c
32c3540c
0a7403e4
0010603c
16c305c3
0ae328bc
11940007
343cd40f
546c100c
07c38d00
6ebc2386
60260a7c
000d033c
03a3700c
0006100f
08040f56
0136f016
71c340c3
0ae3acbc
238607c3
0a7c5cbc
503c80c3
04c30010
28bc15c3
60c30ae3
b00f0df2
07c3906c
6ebc2386
60260a7c
000d033c
043c38c3
06c33b9d
0f568076
00000804
fc96f016
71c360c3
5ebc0fc3
40c30ae2
18940007
06bc06c3
30c30ae3
13c30fc3
0ae964bc
0bf240c3
16c30fc3
30bc2fc3
40c30ae6
60d704f2
5c0f4c0c
7ebc0fc3
04c30ae2
0f560496
00000804
0f36f016
b1c380c3
200c62c3
32c3482c
077413e4
202506c3
0ae328bc
3e940007
18c35810
384f244c
287028c3
8006f86c
03b354c3
20060bc3
233c39c3
31c35a1d
0a7e5abc
100031c3
04e42026
20060214
20c36580
ffff101c
0fff111c
273c2183
203c027f
433ce08c
a025212c
680c28c3
51e413c3
9c0fe074
37c325c3
20060073
40252c0f
2ae46085
28c3fb74
6025680c
06c3780f
0ae3bebc
f0760006
08040f56
0136f016
41c350c3
502c200c
13e432c3
04c30774
28bc2025
00070ae3
f00c3194
d00fd40c
106c1470
31c32006
68c30213
1a1d263c
09ac323c
ffff601c
0fff611c
303c3683
2025027f
d88c323c
62c3540c
ee7416e4
202666d2
700c200f
700f6c80
323c500c
d06c100c
00b36f00
133c2006
4025027f
fb7427e4
304f344c
80760006
08040f56
50c37016
0020613c
10f8301c
0000311c
8c0c6c0c
100c063c
41262006
681c301c
0016311c
30c34664
1fc6146f
20066fd2
d42f340f
21c3344f
746c00d3
133c2006
40252b9d
fa7426e4
0e560006
00000804
3f36f016
0077fc96
600cc1c3
080cd33c
3de4642c
01c30815
28bc1dc3
00070ae3
000c54dc
d31c1f86
06dc0200
301c000c
311c10f8
6c0c0000
001c8c0c
20060800
301c4126
311c680c
46640016
1fc600b7
40074097
000ab2dc
a6c3c006
0eb3c037
fff0233c
02f436e4
192026c3
64702057
21e42c20
123c0315
303c0010
4bc3100c
80f79180
100c323c
93849bc3
0010323c
61526c20
13e481c3
83c302f4
54c38006
02b374c3
040c19c3
60d72006
4a1d233c
5abc31c3
14000a7e
05e44026
40060214
50c37c80
921ce980
8025fffc
eb7448e4
080c253c
25e42026
20060214
080c373c
4ac36580
2026aa00
021452e4
40172006
e5806d00
17c325c3
0014463c
14948007
090c363c
303c0bc3
03c33a1d
23c314c3
5abc34c3
31c30a7e
20265400
021425e4
7d8014c3
32c32580
ffff401c
0fff411c
00973483
6b9d303c
e08ca23c
252ca13c
e08c313c
c0256037
700c8057
89746de4
040c1cc3
640f6112
4006246c
80970193
2a1d343c
ffff401c
0fff411c
313c3483
4025027f
f4742de4
800600b3
027f413c
20e44025
0cc3fb74
0ae3bebc
10f8301c
0000311c
8c4c6c0c
20060097
301c4126
311c680c
46640016
04960006
0f56fc76
00000804
3f36f016
0037fe96
b2c3d1c3
682c43c3
081534e4
14c302c3
0ae328bc
44dc0007
1dc30009
4017640c
6d00480c
43e4a4c3
a3c302f4
a31c1f86
66dc0200
301c0008
311c10f8
6c0c0000
001c8c0c
20060800
301c4126
311c67f8
46640016
1fc6c0c3
20071cc3
80067154
94c374c3
2dc30893
233c680c
34e4fff0
24c302f4
00173120
3dc3a06c
c0170c6c
83c3780c
28e481a4
823c0315
313c0010
7580100c
323c6077
c180100c
02b3a006
2006180c
233c6057
31c35a1d
0a7e5abc
40261c00
021407e4
79c34006
70c37c80
938492c3
a025df85
eb7458e4
201c37c3
211cffff
32830fff
363c6cc3
373c4b9d
793ce08c
993c21ac
8025e08c
bc744ae4
280c2bc3
486c4811
00f36006
663c6cc3
623c3a1d
6025027f
f915a3e4
000600b3
027f023c
31e46025
0bc3fb74
0ae3bebc
10f8301c
0000311c
8c4c6c0c
20060cc3
301c4126
311c67f8
46640016
02960006
0f56fc76
00000804
50c3f016
01c371c3
0ae306bc
c027dc0c
23860ef4
0a7c6ebc
363c40c3
7c6501c7
2e0005c3
0ae964bc
03d307d2
202605c3
0ae56cbc
9fe58026
05c30293
febc15c3
00070ae9
05c31194
1ebc17c3
1fe70ae5
05c30754
25c317c3
0ae630bc
802505f2
ecf48367
0f560006
00000804
fc96f016
71c360c3
5ebc0fc3
40c30ae2
14940007
06bc06c3
30c30ae3
13c30fc3
0ae964bc
07f240c3
16c30fc3
30bc27c3
40c30ae6
7ebc0fc3
04c30ae2
0f560496
00000804
3f36f016
0077fa96
a2c3d1c3
640c6037
8c00000c
34e4682c
02c30815
28bc14c3
00070ae3
0009f4dc
431c1f86
a6dc0200
301c0009
311c10f8
6c0c0000
001c8c0c
20060800
301c4126
311c67e0
46640016
1fc600b7
60076097
000852dc
700c4dc3
c057c3c3
c084180c
02120017
20970137
b084b1c3
00048f5c
00a7bf5c
94c38006
2dc308b3
233c680c
38e4fff0
28c302f4
212008c3
ac6c6057
186c6dc3
eca06c0c
031527e4
0010723c
100c313c
60f77580
100c323c
a006c180
180c02b3
60d72006
5a1d233c
5abc31c3
10000a7e
04e44026
40060214
708049c3
92c340c3
df859384
57e4a025
34c3eb74
ffff201c
0fff211c
c1573283
027f363c
343cc177
493ce08c
993c21ac
821ce08c
8ce40001
2ac3bb74
8811280c
8117686c
60174e00
6bc30113
0004b21c
623cd80c
6025027f
f8f43ce4
800600b3
027f423c
31e46025
0ac3fb74
0ae3bebc
10f8301c
0000311c
8c4c6c0c
20060097
301c4126
311c67e0
46640016
06960006
0f56fc76
00000804
40c3f016
acbc61c3
a0060ae3
208604c3
92bc24c3
70c30ae4
12940007
363c506c
280ce08c
680f31a3
6025700c
a025700f
0354a107
fd73c412
bebc04c3
07c30ae3
08040f56
0336f016
81c360c3
200c72c3
20c3082c
087412e4
202507c3
0ae328bc
000740c3
b84c5894
0f94a027
184f0006
18c306c3
86bc27c3
40c30aed
b84fbc4f
bebc07c3
08f30ae3
186c3c10
780c5c6c
05946027
18e4200c
02130435
01d367d2
74a058c3
027f323c
823c0073
0026027f
1c0f1c4f
31c310c3
20060513
780c3c4f
600c7c0f
433c38a4
501cf88c
511cffff
35830fff
027f323c
01d32026
1a1d303c
433c6e20
501cf88c
511cffff
35830fff
027f323c
780c2025
15e453c3
fb93f074
023c0006
6025027f
fb7439e4
bebc07c3
80060ae3
c07604c3
08040f56
0136f016
71c350c3
200c62c3
20c3082c
087412e4
202506c3
0ae328bc
000740c3
744c6694
17946027
6027740c
746c05d4
37e46c0c
60061014
05c3744f
26c317c3
0aed1abc
e02640c3
f44ff84f
bebc06c3
09b30ae3
00061810
346c184f
744c586c
2b946007
7c00040c
e08c433c
ffff701c
0fff711c
323c3783
0026027f
713c01d3
73800a1d
e08c433c
ffff701c
0fff711c
323c3783
0025027f
73c3740c
f07407e4
382c88d2
03e431c3
00250415
027f423c
6025740c
02b3780f
180f0026
423c140c
00270040
a40c0694
680f7ea0
013324c3
24c3e80f
00b30026
723ce006
0025027f
fb7408e4
bebc06c3
80060ae3
807604c3
08040f56
40c31016
4006000c
03f210c3
40250373
051520e4
333c706c
7ad22a1d
033c706c
123c2a1d
303c01c7
6cf20014
67a0201c
0016211c
00f4303c
3a1d423c
04322600
01c37ad2
08040856
00073016
303c1154
3083fff0
23c36df2
343c8026
03e4200d
440f0494
00b30026
43874025
0006f794
08040c56
0736f016
50c3ff96
72c361c3
0ae3acbc
ffe0373c
67c71fa6
780845b4
0000801c
049465a7
801cc025
05c30001
0ae3acbc
6394a01c
0016a11c
1474901c
0000911c
e4670533
40370ed4
600c0ac3
31c32d22
0002341c
5c0563d2
2f5c4037
20640001
200c09c3
66028006
045432e4
88078025
47e4fb94
05c31215
25c317c3
0ae9aebc
10940007
14c305c3
86bc25c3
0af20aed
5808c025
d6944007
03c3740c
145163d2
01960006
0f56e076
00000804
fc967016
51c340c3
14c30fc3
b0bc4206
04c308cb
420615c3
08cbb0bc
1fc305c3
b0bc4206
049608cb
08040e56
3f36f016
c0c3f696
40b7a1c3
400cd3c3
2d00640c
01fe131c
32e40fd4
32c302f4
00ff331c
0cc309d4
40971ac3
42bc3dc3
b0c30aec
0f3c0cb3
20250180
0aea40bc
0007b0c3
1cc35d94
2077240c
480c2ac3
60256500
40f761b7
100c0d3c
90c30177
07d36bc3
646c1cc3
6a1d333c
62576137
ad004157
86a48dc3
706c4ac3
ec0009c3
04d38006
20060117
31c35c0c
0a7e5abc
203730c3
4c80340c
23e42026
20060214
64000017
20260a00
021402e4
65802006
20c3e085
ffff101c
0fff111c
253c2183
203c027f
433ce08c
821c212c
40d70001
83e432c3
940fd874
921cc025
8057fffc
60e404c3
4f3cc074
04c30180
0ae3bebc
209704c3
0aee90bc
7ebc04c3
0bc30ae2
fc760a96
08040f56
3f36f016
b0c3f896
4077c1c3
331c93c3
12d401ff
1bc3440c
32e4640c
32c302f4
00ff331c
0bc309d4
40571cc3
42bc39c3
a0c30aeb
0f3c0c33
19c30100
0aea40bc
0007a0c3
9f5c5994
1bc30087
20b7240c
085340c3
84a489c3
780c6cc3
02f483e4
1bc383c3
333c646c
60f74a1d
100c343c
ed0041d7
ac703cc3
65c3a006
00d704d3
3dc32006
5a1d233c
5abc31c3
30c30a7e
1c0c2037
20264c00
021423e4
00172006
0b006400
02e42026
20060214
20c36580
ffff101c
0fff111c
273c2183
203c027f
633ce08c
a025212c
da7458e4
39e47600
dc0f0215
20978025
42e421c3
4f3cbc74
04c30100
0ae3bebc
205704c3
0aee90bc
7ebc04c3
0ac30ae2
fc760896
08040f56
0136f016
52c341c3
e44cc04c
500c200c
60256500
01ff331c
21e40cd4
21c302f4
0100231c
14c306d4
42bc25c3
00b30aeb
25c314c3
0aef2abc
4006740c
07f432e4
363c6703
33c40b0d
f88c233c
8076544f
08040f56
0336f016
50c3fc96
82c391c3
0fc3e40c
8abc15c3
40c30ae3
62940007
173c0fc3
f4bcfff0
40060ae3
0800211c
73e432c3
0fc30735
2fc318c3
0aefaabc
0fc300f3
2fc318c3
a6bc37c3
40c30aee
45940007
0fc3e025
f4bc17c3
05c30ae3
01c7173c
1abc25c3
40c30ae4
37940007
19c30fc3
37c32fc3
0aef2abc
000740c3
05c32e94
25c31fc3
0ae698bc
000780c3
05c32594
5abc18c3
1fe70ae5
0fc31994
6cbc2026
0fc30ae5
62bc17c3
40c30ae4
15940007
1fc305c3
7abc25c3
00d30ae6
19c305c3
30bc25c3
40c30ae6
05c308f2
42bc19c3
1fe70ae5
48c3f494
7ebc0fc3
04c30ae2
c0760496
08040f56
3f36f016
b0c3f796
40102077
080c3a3c
0010433c
01400f3c
40bc14c3
d0c30aea
84dc0007
81770009
c01c5dc3
10730004
180c353c
8c802217
100c653c
686c2bc3
5a1d333c
200603c3
31c323c3
0a7e5abc
21c330c3
0380f00c
03e42026
20060214
30c34500
ffff101c
0fff111c
700f3183
e08c303c
21ac423c
686c2bc3
60f76f01
3c846217
253c6137
40b70010
72c385c3
63c3e212
1bc305f3
0f81646c
40d72006
5abc31c3
91c30a7e
5180780c
20372026
031424e4
80378006
20268800
021442e4
40172006
398432c3
10006580
04e42026
20060214
45803984
401c30c3
411cffff
34830fff
027f363c
e08c303c
21ac423c
821ce085
8ae40001
35e3cf74
62123a84
29804117
640c0273
00265180
021424e4
32c30006
ffff401c
0fff411c
313c3483
323c027f
403ce08c
800721ac
c21ced94
a0970008
d3dc5ae4
4f3cfff7
04c30140
0ae3bebc
205704c3
0aee90bc
7ebc04c3
0dc30ae2
fc760996
08040f56
40c37016
400c51c3
080c323c
01fe331c
4fe706d4
68bc04d4
00b30aea
15c304c3
0af048bc
d44fc006
08040e56
3f36f016
b0c3fa96
d2c32077
00800f3c
280c2bc3
0aea40bc
0007c0c3
5bc37594
60b7740c
0137144c
fff0a33c
100c8a3c
1cc34cc3
343c0a93
713c208c
2bc3e1ac
58c3686c
443c6e81
17c3e1ac
67c3e4f2
3e358047
17c304c3
5555201c
0555211c
5abc6006
603c0a7e
613ce08c
513c232c
16c4e08c
22f24026
35c421c3
92a493c3
60264720
21e46037
600603b4
09c36037
a01762a0
0a006ea0
02e48026
80060214
71806f80
2026a080
021450e4
39842006
05c38580
406614c3
e0bc6006
c3000a7d
14c305c3
60064066
0a7e22bc
615740c3
cee158c3
ffffa21c
fffc821c
0000a31c
2dc3ab15
880f42d2
6ad26057
00804f3c
bebc04c3
04c30ae3
90bc2057
0f3c0aee
7ebc0080
0cc30ae2
fc760696
08040f56
0336f016
90c3fc96
72c351c3
200783c3
12c30cd4
0ae35abc
38c340c3
3c546007
acbc08c3
07130ae3
5ebc0fc3
40c30ae2
32940007
69d238c3
15c309c3
1abc2fc3
40c30ae4
25940007
17c309c3
0ae35abc
000740c3
a3671e94
05c30af4
5cbc2386
30c30a7c
13c307c3
0ae3f4bc
238605c3
0a7c6ebc
04d210c3
d4bc07c3
07c30ae3
0ae3bebc
65d238c3
18c30fc3
0aee90bc
7ebc0fc3
04c30ae2
c0760496
08040f56
0336f016
50c3fc96
92c361c3
5ebc0fc3
40c30ae2
2c940007
06bc06c3
80c30ae3
18c305c3
35c32fc3
0af194bc
000740c3
0fc31c94
2fc319c3
0aefaabc
000740c3
05c31494
25c31fc3
0ae5d2bc
0df240c3
16c305c3
0ae51ebc
07541fe7
16c305c3
30bc25c3
fbb30ae6
7ebc0fc3
04c30ae2
c0760496
08040f56
0336f016
50c3fc96
82c361c3
5ebc0fc3
40c30ae2
2f940007
06bc06c3
90c30ae3
19c305c3
35c32fc3
0af194bc
000740c3
831c1f94
09540001
18c30fc3
aebc2fc3
40c30ae9
14940007
1fc305c3
d2bc25c3
40c30ae5
05c30df2
1ebc16c3
1fe70ae5
05c30754
25c316c3
0ae630bc
0fc3fb53
0ae27ebc
049604c3
0f56c076
00000804
fc96f016
71c330c3
13c30fc3
0ae38abc
40c350c3
02d30ed2
4c0960d7
0fc35ea1
2fc32106
94bc6006
40c30af1
a02508f2
93f28017
15c307c3
0ae396bc
7ebc0fc3
04c30ae2
0f560496
00000804
fc963016
0fc330c3
8abc13c3
50c30ae3
a0060ed2
60d70233
533c6c0c
0fc309cb
2fc32106
94bc6006
03f20af1
74f26017
7ebc0fc3
05c30ae2
0c560496
00000804
0136f016
40c3f896
82c351c3
63f2600c
007301c3
66f2640c
12bc18c3
40c30ae5
7f3c1013
07c30100
8abc14c3
40c30ae3
77940007
15c30fc3
0ae38abc
000740c3
00b76d94
07c301b7
0aee00bc
0fc350c3
0aee00bc
60c370c3
02f405e4
c00765c3
0f3c14f4
16c30100
600620c3
0af194bc
000740c3
0fc34f94
2fc316c3
94bc34c3
40c30af1
46940007
0b5456e4
01000f3c
20c33720
94bc6006
40c30af1
3a940007
2a5476e4
3f200fc3
60062fc3
0af194bc
000740c3
04132f94
1fc307c3
0ae51ebc
05940027
1fc307c3
0aee90bc
17c30fc3
30bc2fc3
40c30ae6
1c940007
00bc0fc3
30c30aee
13c30fc3
34c32fc3
0af194bc
04d240c3
7f3c01f3
60170100
dd946007
16c307c3
92bc28c3
40c30ae4
38c303f2
0f3c0c4f
7ebc0100
0fc30ae2
0ae27ebc
089604c3
0f568076
00000804
3f36f016
60c3fb96
a2c371c3
bfa683c3
c2dc2007
20270008
780c0354
18c36df2
400623d2
3ac3440f
7f546007
1ac306c3
0ae35abc
01c30493
01001f3c
0aee24bc
16940027
4bd228c3
00833f5c
303c0323
586cfff0
3083080c
640f18c3
40072ac3
06c36454
60062117
0af194bc
e0670113
06c30894
28c31ac3
0af10cbc
0ad350c3
380c0fc3
0aea40bc
000750c3
780c4f94
184c6037
7fe500b7
45c36137
d5c315c3
343c05f3
913c208c
786ce1ac
333c1bc3
443c1a1d
19c3e1ac
0594d9e4
0000c01c
17b474e4
19c304c3
600627c3
0a7de0bc
2006c0c3
31c327c3
0a7e5abc
502031c3
24e42026
200602b4
61a009c3
2ca042c3
2bc360d7
2b9dc33c
7fe56117
bf5c6137
b31c0084
ce150000
02d208c3
1ac3800f
0fc328d2
0ae3bebc
1ac30fc3
0aee90bc
7ebc0fc3
00530ae2
05c3a006
fc760596
08040f56
400632c3
0af33cbc
00000804
0136f016
60c3ff96
400651c3
401c440f
411c63a0
701c0016
711c6398
06c30016
2fc3300c
0af3d6bc
60170af2
602664f2
00b3740f
7c0c8085
f29443e4
80760196
08040f56
3f36f016
d0c3ed96
a2c3c1c3
640c63c3
60079fa6
000b92dc
0ae51ebc
10941fe7
c6d246c3
16c30dc3
0ae35abc
3ac340c3
a2dc6007
0ac3000a
0ae3acbc
bf3c14b3
8f3c03c0
9f3c02c0
400601c0
40774037
18c30bc3
3f3c29c3
a4bc00c0
40c30ae2
24dc0007
09c30009
6cbc2026
0dc30ae5
0ae306bc
0cc370c3
0ae306bc
0dc350c3
12bc1bc3
40c30ae5
6e940007
18c30cc3
0ae512bc
000740c3
bea06794
15c308c3
92bc28c3
40c30ae4
5e940007
15c309c3
92bc29c3
00b70ae4
55940007
89c378c3
07c30573
42bc1bc3
00270ae5
0bc31254
2bc317c3
0ae698bc
000740c3
0f3c4594
18c300c0
7abc20c3
40c30ae6
3c940007
202607c3
600627c3
0af194bc
000740c3
08c33394
28c32026
94bc34c3
40c30af1
0007bfe5
a0072994
2dc3d515
3cc3884c
2ac3ac4c
13544007
1f3c0ac3
90bc00c0
2ac30aee
03c3680c
34c368d2
333c3503
33c40b0d
f88c033c
0c4f3ac3
06c3ccd2
03c01f3c
0aee90bc
62f2780c
984f43c3
00538006
0f3c8097
7ebc03c0
0f3c0ae2
7ebc02c0
0f3c0ae2
7ebc01c0
0f3c0ae2
7ebc00c0
04c30ae2
fc761396
08040f56
0336f016
60c3f696
82c351c3
01807f3c
00809f3c
40374006
07c34077
32c319c3
0ae2a4bc
000740c3
06c33394
27c315c3
0af2a6bc
000740c3
06c32394
1ebc15c3
1fe70ae5
06c30c94
29c317c3
febc34c3
40c30af3
800705c3
01531394
17c305c3
34c329c3
0af3febc
0af240c3
19c306c3
aabc28c3
40c30aef
38c34006
0f3c4c4f
7ebc0180
0f3c0ae2
7ebc0080
04c30ae2
c0760a96
08040f56
50c33016
640c41c3
0387133c
0ae964bc
07f230c3
14c305c3
febc25c3
30c30af3
0c5603c3
00000804
0136f016
70c3fc96
82c351c3
5ebc0fc3
40c30ae2
1d940007
15c307c3
3fc324c3
0af3febc
000740c3
60971194
21c3344c
085432e4
1fc305c3
7abc28c3
40c30ae6
0fc300b3
90bc18c3
0fc30aee
0ae27ebc
049604c3
0f568076
00000804
0136f016
60c3fc96
82c371c3
5ebc0fc3
40c30ae2
10940007
1fc306c3
0af0f6bc
07f240c3
17c30fc3
26bc28c3
40c30af5
7ebc0fc3
04c30ae2
80760496
08040f56
0336f016
60c3fc96
82c371c3
0fc393c3
0ae25ebc
000740c3
06c31194
2fc317c3
0aefaabc
07f240c3
18c30fc3
26bc29c3
40c30af5
7ebc0fc3
04c30ae2
c0760496
08040f56
3f36f016
fdc8f21c
207780c3
6037b2c3
06bc01c3
c01c0ae3
00e70002
c01c0cf4
04870003
c01c08f4
031c0005
03d4008c
0004c01c
02800f3c
0ae25ebc
000740c3
0016b4dc
fff07c3c
233c6026
4177700d
c00d233c
415740b7
3f3c4412
4d000180
c1574137
035352c3
5ebc05c3
40c30ae2
0007a205
a1571254
01170133
0ae27ebc
6117a025
220513c3
56e42137
0f3cf774
7ebc0280
28130ae2
6097c025
61e413c3
5f3ce474
05c32180
0ae25ebc
000740c3
0011e4dc
13242f5c
05c34ef2
12bc1bc3
40c30af5
f4dc0007
a01c0010
a11cdfa8
01b30015
15c30bc3
0aec20bc
000740c3
001024dc
e3c8a01c
0015a11c
02805f3c
1bc308c3
26bc25c3
40c30af5
34dc0007
6206000f
700d233c
01803f3c
05c3cd00
5abc16c3
40c30ae3
54dc0007
50c3000e
21808f3c
16c306c3
0af0f6bc
000740c3
000da4dc
1bc306c3
a66428c3
000740c3
000d24dc
57e4a025
2157ee74
c02561c3
200c263c
01803f3c
e117ad00
02809f3c
07c302b3
25c319c3
0aefaabc
000740c3
000ba4dc
1bc305c3
a66428c3
a20540c3
0007e205
000b04dc
4097c025
63e432c3
8f3ce974
08c32280
0ae25ebc
000740c3
000a24dc
202608c3
0ae56cbc
640c2057
fff0133c
d4c320f7
64c374c3
0001901c
007354c3
080cdd3c
ffff921c
4ef229c3
13c360d7
52543fe7
686c4057
d33c20d7
3fe51a1d
901c20f7
2d3c001c
32c30ecb
63f235a3
fcf353c3
1094a027
08c34ff2
f6bc18c3
00070af0
08c36094
2f3c1bc3
a6642180
d7540007
c0250b13
67201cc3
300d323c
a04673a3
cd946ce4
08c3a006
f6bc18c3
00070af0
08c34894
2f3c1bc3
a6642180
41940007
5ce4a025
373cf174
08c3200c
01802f3c
28c32980
0aefaabc
33940007
1bc308c3
21802f3c
0007a664
70c32c94
a02660c3
a047f4d3
c0072b94
59c329f4
22808f3c
21809f3c
0280cf3c
18c308c3
0af0f6bc
17940007
1bc308c3
a66429c3
11940007
37c3e112
32834097
08c36ed2
28c31cc3
0aefaabc
08c306f2
29c31bc3
03d2a664
013340c3
56e4a025
0f3ce074
20172280
0aee90bc
22800f3c
0ae27ebc
21800f3c
0ae27ebc
02800f3c
0ae27ebc
01170193
0ae27ebc
21c32157
41774025
13c36117
21372205
32c34157
32e44097
04c3f174
0238f21c
0f56fc76
00000804
3f36f016
fdd4f21c
207780c3
603792c3
06bc01c3
20460ae3
00e720f7
60660cf4
048760f7
40a608f4
031c40f7
03d4008c
20f72086
02800f3c
0ae25ebc
000740c3
001ad4dc
72c340d7
6026ffe5
700d233c
20d74177
100d233c
415740b7
3f3c4412
4d000180
c1574137
035352c3
5ebc05c3
40c30ae2
0007a205
a1571254
01170133
0ae27ebc
4117a025
620532c3
56e46137
0f3cf774
7ebc0280
30130ae2
4097c025
63e432c3
1f5ce474
200712c4
09c31994
22801f3c
0ae724bc
000740c3
0015a4dc
4c0c39c3
080c323c
01fe331c
231c24d4
21d400ff
ce9cb01c
0015b11c
1f3c0413
2f5c2280
32c312c4
09946027
d4bc09c3
b01c0ae8
b11cd1b8
02330015
88bc09c3
40c30ae9
54dc0007
b01c0013
b11ce440
00b30015
d09cb01c
0015b11c
21805f3c
5ebc05c3
40c30ae2
34dc0007
1f5c0012
200712c4
05c31194
eabc19c3
40c30aeb
34dc0007
08c30011
29c315c3
02803f3c
0af574bc
05c30173
6cbc2026
08c30ae5
2f3c19c3
26bc0280
40c30af5
d4dc0007
6206000f
700d233c
01803f3c
0f3ccd00
16c30280
0ae35abc
000740c3
000ee4dc
06c350c3
f6bc16c3
40c30af0
54dc0007
06c3000e
2f5c19c3
b6641144
40c303d2
a0251b93
ee7457e4
63c36157
263cc025
3f3c200c
ad000180
8f3ce117
02d30280
18c307c3
aabc25c3
40c30aef
54dc0007
05c3000c
2f5c19c3
b6641144
a20540c3
0007e205
000ba4dc
2097c025
62e421c3
2057e874
d33c640c
c006fff0
76c386c3
0001c01c
af3c56c3
00532180
c21cc112
2cc3ffff
d31c4df2
5c54ffff
646c2057
633c2dc3
d21c2a1d
c01cffff
263c001c
32c30ecb
63f235a3
fd3353c3
1494a027
12944007
1ac30ac3
0af0f6bc
000740c3
000844dc
19c30ac3
11442f5c
40c3b664
d5540007
e0250f53
67a020d7
300d323c
a04683a3
cb9471e4
0ac3a006
f6bc1ac3
40c30af0
69940007
19c30ac3
11442f5c
40c3b664
61940007
60d7a025
51e413c3
383ced74
0ac3200c
01802f3c
2ac32980
0aefaabc
000740c3
0ac35094
2f5c19c3
b6641144
000740c3
80c34894
a02670c3
a047f3d3
e0073194
5cc32ff4
21806f3c
0280af3c
16c306c3
0af0f6bc
000740c3
06c33494
2f5c19c3
b6641144
000740c3
883c2c94
38c3080c
32834097
11546007
1ac306c3
aabc26c3
40c30aef
1d940007
19c306c3
11442f5c
40c3b664
15940007
57e4a025
1f5cd874
29f212c4
21800f3c
2f5c19c3
b6641144
07f240c3
21800f3c
90bc2017
80060aee
21800f3c
0ae27ebc
02800f3c
0ae27ebc
01170193
0ae27ebc
32c34157
61776025
21c32117
41374205
13c36157
13e46097
04c3f174
022cf21c
0f56fc76
00000804
1f36f016
50c3de96
c2c361c3
6027644c
001872dc
6007640c
001832dc
07807f3c
06808f3c
03803f3c
3f3c6037
60770280
18c307c3
05802f3c
04803f3c
0ae2a4bc
000740c3
001834dc
00770037
01800f3c
00801f3c
34c324c3
0ae2a4bc
000740c3
001754dc
16c305c3
26bc27c3
40c30af5
54dc0007
06c30013
5abc18c3
40c30ae3
d4dc0007
67970012
10f46007
6c0c6857
0001341c
66976bf2
08f46007
6c0c6757
0001341c
a2dc6007
9f3c0011
09c30780
05801f3c
0ae35abc
000740c3
001104dc
06807f3c
04805f3c
15c307c3
0ae35abc
000740c3
001044dc
03800f3c
6cbc2026
4f3c0ae5
04c30080
6cbc2026
a5c30ae5
01808f3c
54c3b7c3
073379c3
60076397
001117dc
6c0c6457
0001341c
a2dc6007
00f30010
6c0c6357
0001341c
15546007
03800f3c
20c31bc3
0ae67abc
000740c3
000d64dc
02800f3c
20c317c3
0ae698bc
000740c3
000cc4dc
03800f3c
94bc10c3
40c30ae5
34dc0007
0f3c000c
10c30280
0ae594bc
000740c3
000ba4dc
60076597
665742f4
341c6c0c
60070001
0f3c3c94
10c30580
0ae594bc
000740c3
14f3b854
60076197
000cc7dc
6c0c6257
0001341c
52dc6007
00f3000c
6c0c6157
0001341c
13546007
1bc308c3
7abc28c3
40c30ae6
d4dc0007
05c30008
25c317c3
0ae698bc
000740c3
000844dc
18c308c3
0ae594bc
000740c3
05c37c94
94bc15c3
40c30ae5
75940007
60076497
0009f7dc
6c0c6557
0001341c
84dc6007
0ac30009
94bc1ac3
40c30ae5
bd540007
04c30c53
24c31ac3
0ae698bc
000740c3
0f3c5a94
18c30380
98bc20c3
40c30ae6
51940007
02800f3c
20c315c3
0ac302d3
2ac314c3
0ae698bc
000740c3
08c34494
03801f3c
98bc28c3
40c30ae6
3b940007
1f3c05c3
25c30280
0ae698bc
000740c3
65973294
74dc6007
0f3cfff7
20260480
0ae55abc
26940007
05c30133
25c316c3
0ae67abc
04d240c3
5f3c03d3
05c30180
5abc2006
1fe70ae5
0113f154
16c305c3
98bc25c3
40c30ae6
05c30ef2
1ebc16c3
1fe70ae5
05c3f494
90bc1cc3
80060aee
9fa60053
07800f3c
0ae27ebc
06800f3c
0ae27ebc
05800f3c
0ae27ebc
04800f3c
0ae27ebc
03800f3c
0ae27ebc
02800f3c
0ae27ebc
01800f3c
0ae27ebc
00800f3c
0ae27ebc
9fa602f3
629702b3
76dc6007
e1f3ffef
60076097
fff3c6dc
4f3cea53
04c30580
42bc1ac3
1fe70ae5
fff6b4dc
04c3eff3
f8762296
08040f56
3f36f016
d0c3e596
40b7b1c3
6007640c
000e57dc
6c0c646c
0001341c
60079fa6
000fc2dc
0bc31b73
5abc17c3
40c30ae3
b4dc0007
0dc3000b
25c31bc3
0af526bc
000740c3
000b24dc
19c307c3
0ae35abc
000740c3
000aa4dc
18c305c3
0ae35abc
40c350c3
14dc0007
06c3000a
6cbc2026
a5c30ae5
5cc379c3
61d70353
10f46007
6c0c6297
0001341c
05c36bd2
05c01f3c
98bc25c3
40c30ae6
74dc0007
05c30008
94bc15c3
40c30ae5
7f940007
600763d7
649727f4
341c6c0c
60070001
07c32194
94bc17c3
40c30ae5
d8540007
60d70dd3
0ff46007
6c0c6197
0001341c
06c36ad2
05c01f3c
98bc26c3
40c30ae6
5d940007
16c306c3
0ae594bc
000740c3
62d75694
47dc6007
63970008
341c6c0c
60070001
08c37d94
94bc18c3
40c30ae5
d8540007
07c30893
27c318c3
0ae698bc
000740c3
05c33c94
25c316c3
08c30193
28c317c3
0ae698bc
000740c3
06c33094
26c315c3
0ae698bc
000740c3
63d72894
a21c67d2
a31c0001
a3f41000
0f3c03f3
202602c0
0ae55abc
18940007
c84c2dc3
00c05f3c
05c30113
25c31bc3
0ae67abc
0df240c3
60276157
05c3f754
90bc2097
60970aee
8006cc4f
9fa60053
05c00f3c
0ae27ebc
04c00f3c
0ae27ebc
03c00f3c
0ae27ebc
02c00f3c
0ae27ebc
01c00f3c
0ae27ebc
00c00f3c
0ae27ebc
7f3c0413
5f3c05c0
9f3c04c0
8f3c03c0
cf3c02c0
cf5c01c0
6f3c0007
c07700c0
15c307c3
38c329c3
0ae2a4bc
09f240c3
07c3e1f3
42bc18c3
1fe70ae5
f2538794
1b9604c3
0f56fc76
00000804
50c3f016
62c341c3
6027644c
640c0d54
60076bd2
646c0bf4
341c6c0c
66d20001
0afaa6bc
1fa60113
05c300d3
26c314c3
0af8fcbc
08040f56
0336f016
70c3f596
52c381c3
401c93c3
411c10f8
900c0000
4664906c
3f5c00b7
43c30041
65546007
9fa6744c
61546027
684c28c3
2d946027
01c06f3c
5ebc06c3
40c30ae2
55940007
15c307c3
b8bc26c3
40c30afb
7f3c08f2
07c300c0
0ae25ebc
03d240c3
025306c3
17c308c3
0ae512bc
08f240c3
17c306c3
39c325c3
0afbd4bc
06c340c3
0ae27ebc
7ebc07c3
06330ae2
bcbc05c3
00270ae6
05c32454
0ae70cbc
05c305f2
0ae6e2bc
740c0112
32e44006
40060df4
6c0c746c
0001341c
402662f2
0016123c
2f5c2077
40270021
09d20254
07c30037
25c318c3
28bc39c3
01130af7
07c30037
25c318c3
96bc39c3
40c30af5
0b9604c3
0f56c076
00000804
1f36f016
90c3f496
c2c3a1c3
680f6006
202601c3
0ae55abc
9fa670c3
75940027
02008f3c
19c308c3
0ae38abc
000740c3
08c36c94
28c317c3
0aed1abc
000740c3
0fc36094
8abc18c3
40c30ae3
59940007
00bc0fc3
b0c30aee
1bc30fc3
34c32fc3
0af194bc
000740c3
6f3c4994
06c30100
0ae25ebc
000740c3
0ac34194
29c31fc3
d4bc36c3
a0c30afb
33940007
17c306c3
0ae55abc
28540007
18c306c3
0ae542bc
22540007
78c357c3
06c30213
26c319c3
0af554bc
000740c3
06c31d94
5abc2026
00070ae5
a0251754
07f4b5e4
17c306c3
0ae542bc
ea940007
01000f3c
02001f3c
0ae542bc
602606f2
680f2cc3
00538006
0f3c4ac3
7ebc0100
0fc30ae2
0ae27ebc
02000f3c
0ae27ebc
0c9604c3
0f56f876
00000804
1f36f016
80c3fb96
92c3b1c3
680f6006
fff0313c
331c9fa6
47b400ff
63a0601c
0016611c
639c401c
0016411c
380c08c3
0ae55abc
402606f2
4c0f39c3
06b340c3
700cc085
f39463e4
0100af3c
1ac308c3
0af3dcbc
000740c3
61172894
25546027
5ebc0fc3
40c30ae2
1f940007
c63c50c3
6ac3c000
0fc30213
133c3cc3
6cbc5a1d
08c30ae5
26c31fc3
0afc52bc
61170af2
a02568d2
f0745be4
39c34026
00534c0f
0fc340c3
0ae27ebc
059604c3
0f56f876
00000804
50c33016
1f540007
0007006c
740c1954
100c133c
0b06b8bc
10f8301c
0000311c
8c4c6c0c
2006146c
301c4126
311c6850
46640016
746f6006
742f740f
6006744f
740f744f
08040c56
ff52001c
00000804
ff52001c
00000804
00000804
01c330c3
023513e4
080403c3
2301201c
6745211c
201c406f
211cab89
408fefcd
dcfe201c
98ba211c
201c40af
211c5476
40cf1032
400f4006
404f402f
00000804
6500402c
32e4602f
604c0434
604f6025
00000804
0336f016
009050c3
80ccc0ac
006c60ec
34c34c00
38833603
09803403
06bc2066
70c30b06
5080350c
380336c3
30c30383
09803603
06bc20e6
40c30b06
5880352c
380337c3
38033083
21660980
0b0606bc
38c360c3
4c00154c
370334c3
37033683
22660980
0b0606bc
356c80c3
36c35c80
30833403
09803403
06bc2066
70c30b06
5180758c
360338c3
36033783
20e60980
0b0606bc
35ac40c3
37c35880
30833803
09803803
06bc2166
60c30b06
15cc38c3
34c34c00
36833703
09803703
06bc2266
80c30b06
5c8035ec
340336c3
34033083
20660980
0b0606bc
760c70c3
38c35180
37833603
09803603
06bc20e6
40c30b06
5880362c
380337c3
38033083
21660980
0b0606bc
38c360c3
4c00164c
370334c3
37033683
22660980
0b0606bc
366c80c3
36c35c80
30833403
09803403
06bc2066
70c30b06
5180768c
360338c3
36033783
20e60980
0b0606bc
36ac90c3
37c35880
30833803
09803803
06bc2166
40c30b06
16cc38c3
39c34c00
34833703
09803703
06bc2266
60c30b06
7d0054ec
7999001c
5a82011c
34c32c00
368339a3
298324c3
058032a3
06bc2066
70c30b06
556c19c3
001c6500
011c7999
2c005a82
34a336c3
26c33783
32a32483
20a60580
0b0606bc
35ec80c3
201c7080
211c7999
2d005a82
36a337c3
27c33083
32a32683
21260580
0b0606bc
166c40c3
201c7800
211c7999
2d005a82
37a338c3
28c33483
32a32783
21a60580
0b0606bc
350c60c3
201c7c80
211c7999
2d005a82
38a334c3
24c33083
32a32883
20660580
0b0606bc
08c370c3
6080358c
7999201c
5a82211c
36c32d00
378334a3
248326c3
058032a3
06bc20a6
80c30b06
7000160c
7999201c
5a82211c
37c32d00
388336a3
268327c3
058032a3
06bc2126
40c30b06
7800168c
7999201c
5a82211c
38c32d00
348337a3
278328c3
058032a3
06bc21a6
60c30b06
7c80352c
7999201c
5a82211c
34c32d00
308338a3
288324c3
058032a3
06bc2066
70c30b06
35ac08c3
201c6080
211c7999
2d005a82
34a336c3
26c33783
32a32483
20a60580
0b0606bc
162c80c3
201c7000
211c7999
2d005a82
36a337c3
27c33883
32a32683
21260580
0b0606bc
16ac40c3
201c7800
211c7999
2d005a82
37a338c3
28c33483
32a32783
21a60580
0b0606bc
354c60c3
201c7c80
211c7999
2d005a82
38a334c3
24c33083
32a32883
20660580
0b0606bc
08c370c3
608035cc
7999201c
5a82211c
36c32d00
378334a3
248326c3
058032a3
06bc20a6
80c30b06
7000164c
7999201c
5a82211c
37c32d00
388336a3
268327c3
058032a3
06bc2126
90c30b06
780016cc
7999201c
5a82211c
38c32d00
398337a3
278328c3
058032a3
06bc21a6
40c30b06
7c8034ec
eba1001c
6ed9011c
39c34c00
34033803
20660980
0b0606bc
28c360c3
680015ec
eba1101c
6ed9111c
34c34c80
36033903
21260980
0b0606bc
29c370c3
6800156c
eba1101c
6ed9111c
36c34c80
37033403
21660980
0b0606bc
566c80c3
001c7100
011ceba1
4c006ed9
360337c3
09803803
06bc21e6
40c30b06
7880352c
eba1001c
6ed9011c
38c34c00
34033703
20660980
0b0606bc
562c60c3
001c7d00
011ceba1
4c006ed9
380334c3
09803603
06bc2126
70c30b06
55ac18c3
001c6500
011ceba1
4c006ed9
340336c3
09803703
06bc2166
80c30b06
708036ac
eba1001c
6ed9011c
37c34c00
38033603
21e60980
0b0606bc
350c40c3
001c7880
011ceba1
4c006ed9
370338c3
09803403
06bc2066
60c30b06
7d00560c
eba1001c
6ed9011c
34c34c00
