36033803
21260980
0b0606bc
18c370c3
6500558c
eba1001c
6ed9011c
36c34c00
37033403
21660980
0b0606bc
368c80c3
001c7080
011ceba1
4c006ed9
360337c3
09803803
06bc21e6
40c30b06
7880354c
eba1001c
6ed9011c
38c34c00
34033703
20660980
0b0606bc
564c60c3
001c7d00
011ceba1
4c006ed9
380334c3
09803603
06bc2126
70c30b06
55cc18c3
001c6500
011ceba1
4c006ed9
340336c3
09803703
06bc2166
80c30b06
708036cc
eba1001c
6ed9011c
37c34c00
38033603
21e60980
0b0606bc
6f00746c
748c746f
748f6c00
388474ac
74cc74af
74cf6f80
0f56c076
00000804
50c3f016
603c71c3
200c01c0
0afd84bc
5006740c
602559a1
6707740f
88060d35
20061980
b0bc51a0
940f0891
8ebc05c3
60060afd
540c740f
20061900
4d206706
0891b0bc
133c744c
542c180c
e88c323c
744f6580
35c34312
027e233c
0380063c
408613c3
08cbb0bc
03c0063c
0080153c
b0bc4086
05c308cb
0afd8ebc
153c07c3
420600c0
08cbb0bc
6abc05c3
0f560afd
00000804
0736f016
81c350c3
903c72c3
a01c01c0
03d30040
07c3940c
2e203ac3
0afd64bc
39c360c3
18c30e00
b0bc26c3
740c08cb
940f9980
0a948807
8ebc05c3
05c30afd
84bc14c3
60060afd
8684740f
e007ff20
e076e294
08040f56
01c330c3
023513e4
080403c3
2301201c
6745211c
201c426f
211cab89
428fefcd
dcfe201c
98ba211c
201c42af
211c5476
42cf1032
400f4006
404f402f
00000804
6500402c
32e4602f
604c0434
604f6025
00000804
0336f016
029050c3
82cce2ac
006c626c
101c6c00
111ca478
4c80d76a
370334c3
34033883
20e60980
0b0606bc
c10028c3
7000148c
b756101c
e8c7111c
37c34c80
06c33803
30c30383
09803703
06bc2186
98000b06
7c8034ac
70db001c
2420011c
36c34c00
34833803
09803803
06bc2226
f0000b06
54cc18c3
001c6500
011cceee
4c00c1bd
360334c3
36033783
22c60980
0b0606bc
808487c3
790054ec
0faf001c
f57c011c
37c34c00
38833403
09803403
06bc20e6
18c30b06
550cc400
001c7100
011cc62a
4c004787
370338c3
37033683
21860980
0b0606bc
552c9800
001c7d00
011c4613
4c00a830
380336c3
38033483
22260980
0b0606bc
18c3f000
6500554c
9501001c
fd46011c
34c34c00
37833603
09803603
06bc22c6
87c30b06
556c8084
001c7900
011c98d8
4c006980
340337c3
34033883
20e60980
0b0606bc
c40018c3
7100558c
f7af001c
8b44011c
38c34c00
36833703
09803703
06bc2186
98000b06
7d0055ac
5bb1001c
ffff011c
36c34c00
34833803
09803803
06bc2226
f0000b06
55cc18c3
001c6500
011cd7be
4c00895c
360334c3
36033783
22c60980
0b0606bc
808487c3
790055ec
1122001c
6b90011c
37c34c00
38833403
09803403
06bc20e6
18c30b06
560cc400
001c7100
011c7193
4c00fd98
370338c3
37033683
21860980
0b0606bc
908496c3
7c00162c
438e101c
a679111c
36c34c80
39833803
09803803
06bc2226
29c30b06
08c38800
6080364c
0821001c
49b4011c
39c34c00
34833603
09803603
06bc22c6
f0000b06
7900548c
2562001c
f61e011c
37c34c00
39833403
09803403
06bc20a6
dc000b06
552c19c3
001c6500
011cb340
4c00c040
370336c3
37033483
21260980
0b0606bc
808486c3
710055cc
5a51001c
265e011c
38c34c00
37833603
09803603
06bc21c6
28c30b06
146c8800
101c7c00
111cc7aa
4c80e9b6
380334c3
38033683
22860980
0b0606bc
550cf000
001c7900
011c105d
4c00d62f
340337c3
34033883
20a60980
0b0606bc
18c3dc00
650055ac
1453001c
0244011c
36c34c00
34833703
09803703
06bc2126
86c30b06
564c8084
001c7100
011ce681
4c00d8a1
360338c3
36033783
21c60980
0b0606bc
880028c3
7c0014ec
fbc8101c
e7d3111c
34c34c80
36833803
09803803
06bc2286
f0000b06
7900558c
cde6001c
21e1011c
37c34c00
38833403
09803403
06bc20a6
dc000b06
562c18c3
001c6500
011c07d6
4c00c337
370336c3
37033483
21260980
0b0606bc
808486c3
710054cc
0d87001c
f4d5011c
38c34c00
37833603
09803603
06bc21c6
28c30b06
156c8800
101c7c00
111c14ed
4c80455a
380334c3
38033683
22860980
0b0606bc
560cf000
001c7900
011ce905
4c00a9e3
340337c3
34033883
20a60980
0b0606bc
18c3dc00
650054ac
a3f8001c
fcef011c
36c34c00
34833703
09803703
06bc2126
86c30b06
554c8084
001c7100
011c02d9
4c00676f
360338c3
36033783
21c60980
0b0606bc
908498c3
480349c3
7c0015ec
4c8a101c
8d2a111c
34c34c80
38033683
22860980
0b0606bc
e80029c3
7800150c
3942101c
fffa111c
47036c80
20860e00
0b0606bc
28c39c00
6800156c
f681101c
8771111c
37c34c80
34033903
21660980
0b0606bc
29c3d000
680015cc
6122101c
6d9d111c
34c34c80
36033703
22060980
0b0606bc
808486c3
7c00162c
380c101c
fde5111c
36c34c80
38033403
22e60980
0b0606bc
e80028c3
7000148c
ea44101c
a4be111c
38c34c80
37033603
20860980
0b0606bc
34ec9c00
001c7880
011ccfa9
4c004bde
380337c3
09803403
06bc2166
d0000b06
554c18c3
001c6500
011c4b60
4c00f6bb
370334c3
09803603
06bc2206
86c30b06
55ac8084
001c7d00
011cbc70
4c00bebf
340336c3
09803803
06bc22e6
18c30b06
560ce400
001c7100
011c7ec6
4c00289b
360338c3
09803703
06bc2086
9c000b06
7900546c
27fa001c
eaa1011c
37c34c00
34033803
21660980
0b0606bc
18c3d000
650054cc
3085001c
d4ef011c
34c34c00
36033703
22060980
0b0606bc
808486c3
7d00552c
1d05001c
0488011c
36c34c00
38033403
22e60980
0b0606bc
e40018c3
7100558c
d039001c
d9d4011c
38c34c00
37033603
20860980
0b0606bc
55ec9c00
001c7900
011c99e5
4c00e6db
380337c3
09803403
06bc2166
d0000b06
564c18c3
001c6500
011c7cf8
4c001fa2
370334c3
09803603
06bc2206
86c30b06
54ac8084
001c7d00
011c5665
4c00c4ac
340336c3
09803803
06bc22e6
18c30b06
546ce400
001c7100
011c2244
4c00f429
17c336e3
31c313a3
09803803
06bc20c6
9c000b06
7900554c
ff97001c
432a011c
38e34c00
13a314c3
370331c3
21460980
0b0606bc
28c3d000
6800162c
23a7101c
ab94111c
37e34c80
03a306c3
340330c3
21e60980
0b0606bc
808486c3
7d00550c
a039001c
fc93011c
34e34c00
03a308c3
360330c3
22a60980
0b0606bc
e40018c3
710055ec
59c3001c
655b011c
36e34c00
13a317c3
380331c3
20c60980
0b0606bc
54cc9c00
001c7900
011ccc92
4c008f0c
14c338e3
31c313a3
09803703
06bc2146
d0000b06
15ac28c3
101c6800
111cf47d
4c80ffef
06c337e3
30c303a3
09803403
06bc21e6
86c30b06
548c8084
001c7d00
011c5dd1
4c008584
08c334e3
30c303a3
09803603
06bc22a6
18c30b06
556ce400
001c7100
011c7e4f
4c006fa8
17c336e3
31c313a3
09803803
06bc20c6
9c000b06
7900564c
e6e0001c
fe2c011c
38e34c00
13a314c3
370331c3
21460980
0b0606bc
28c3d000
6800152c
4314101c
a301111c
37e34c80
03a306c3
340330c3
21e60980
0b0606bc
808486c3
7d00560c
11a1001c
4e08011c
34e34c00
03a308c3
360330c3
22a60980
0b0606bc
e40018c3
710054ec
7e82001c
f753011c
36e34c00
13a317c3
380331c3
20c60980
0b0606bc
908497c3
780015cc
f235101c
bd3a111c
38e34c80
13a319c3
370331c3
21460980
0b0606bc
c80029c3
34ac08c3
001c6080
011cd2bb
4c002ad7
16c337e3
31c313a3
09803903
06bc21e6
98000b06
7d00558c
d391001c
eb86011c
39e34c00
13a314c3
360331c3
22a60980
0b0606bc
3984766c
568c766f
6e006100
76ac768f
76af6e00
6f0076cc
c07676cf
08040f56
50c3f016
603c71c3
200c00c0
0b0108bc
5006740c
602559a1
6707740f
88060d35
20061980
b0bc51a0
940f0891
12bc05c3
60060b01
540c740f
20061900
4d206706
0891b0bc
133c744c
542c180c
e88c323c
744f6580
35c34312
027e233c
0380063c
408613c3
08cbb0bc
03c0063c
0080153c
b0bc4086
05c308cb
0b0112bc
153c07c3
420604c0
08cbb0bc
eebc05c3
0f560b00
00000804
0736f016
81c350c3
903c72c3
a01c00c0
03d30040
07c3940c
2e203ac3
0b00e8bc
39c360c3
18c30e00
b0bc26c3
740c08cb
940f9980
0a948807
12bc05c3
05c30b01
08bc14c3
60060b01
8684740f
e007ff20
e076e294
08040f56
0336f016
71c360c3
901c82c3
911c10f8
29c30000
8c0c680c
20060b86
301c44c6
311c68b8
46640016
706650c3
18540007
0b00eebc
16c305c3
a6bc27c3
05c30b05
5cbc18c3
29c30b05
8c4c680c
200605c3
301c44c6
311c68b8
46640016
03c36006
0f56c076
00000804
6ca06406
318d003c
00000804
118d003c
00000804
20c330c3
ff00101c
ff00111c
48322183
00ff101c
00ff111c
033c3183
2206412c
0b0606bc
00000804
70c3f016
523c61c3
8006108c
063c0113
10bc4a1d
073c0b06
80254b9d
f81445e4
08040f56
0136f016
81c370c3
680642c3
a4bc4d20
50c30a7c
07c361c3
24c318c3
0a7cc2bc
05c350a3
16c361a3
0f568076
00000804
0136f016
81c370c3
680642c3
c2bc4d20
50c30a7c
07c361c3
24c318c3
0a7ca4bc
05c350a3
16c361a3
0f568076
00000804
41c33016
0b0610bc
04c350c3
0b0610bc
0c5615c3
00000804
723cf016
51c3188c
c00640c3
140c0153
66bc342c
100f0b06
c025302f
8105a105
f61467e4
08040f56
51c37016
200642c3
00f321c3
d5016101
61613603
40852025
f91414e4
08040e56
ff967016
61c350c3
31c342c3
20c332a3
32c323a3
0003341c
6ff24006
108c243c
0b0686bc
79220193
752213c3
20371303
00011f5c
40253521
f61424e4
0e560196
00000804
600600b3
00df303c
3cf23fe5
00000804
50c37016
12c341c3
02c34006
d12200f3
d52236c3
03a33603
21e44025
0e56f974
00000804
01c330c3
023513e4
080403c3
028630c3
0e546027
04d46027
6ad20206
040600f3
06546047
60870806
001c0354
0804ff53
22542007
20544007
0f540027
03d40027
035307d2
0d540047
16940087
68060213
6206640f
0253680f
640f6806
00936286
640f6806
680f6406
01130006
0080301c
6806640f
001cff33
0804ff53
3f36f016
b0c3cc96
72c351c3
af5c83c3
cf5c07e4
df5c0804
9f5c0824
931c0844
5db40001
39c3c286
c20662f2
57d4d6e4
0000c31c
39c354f4
16946007
06004f3c
eebc04c3
04c30b00
27c315c3
0b05a6bc
18c304c3
a6bc2ac3
04c30b05
0bc01f3c
0b055cbc
0fc302b3
0b1decbc
39940007
15c30fc3
dabc27c3
0fc30b1d
2ac318c3
0b1ddabc
1f3c0fc3
cabc0bc0
80260b1d
0bc05f3c
06008f3c
931c0313
0b940001
15c30fc3
dabc26c3
0fc30b1d
cabc15c3
01530b1d
15c308c3
a6bc26c3
08c30b05
5cbc15c3
80250b05
e8744ce4
1f3c0bc3
2dc30bc0
08cbb0bc
00730006
ff53001c
fc763496
08040f56
0f36f016
50c3cd96
92c381c3
bf5c73c3
af5c0784
200707a4
0009c2dc
92dc6007
00270009
00272754
08d203d4
00471253
00873e54
0008e4dc
0fc30c93
0b00eebc
18c30fc3
a6bc29c3
0fc30b05
5cbc17c3
a0260b05
0fc30173
2bc317c3
0b05a6bc
17c30fc3
0b055cbc
5ae4a025
8006f574
0fc30e93
0b1decbc
000740c3
0fc36e94
29c318c3
0b1ddabc
17c30fc3
0b1dcabc
0fc30173
2bc317c3
0b1ddabc
17c30fc3
0b1dcabc
5ae4a025
0af3f574
bcbc0fc3
40c30b1d
51940007
18c30fc3
aabc29c3
40c30b1d
49940007
17c30fc3
0b1d9abc
a02680c3
12540007
0fc307f3
2bc317c3
0b1daabc
000740c3
0fc33894
9abc17c3
40c30b1d
31940007
5ae4a025
0593ef74
8cbc0fc3
40c30b1d
27940007
18c30fc3
7abc29c3
40c30b1d
1f940007
17c30fc3
0b1d6abc
a02680c3
10540007
0fc302b3
2bc317c3
0b1d7abc
0ff240c3
17c30fc3
0b1d6abc
09f240c3
5ae4a025
0093f174
ff53401c
48c30053
339604c3
0f56f076
00000804
3f36f016
0137c696
d2c320f7
119760b7
202603f2
121731b7
0dc01f3c
0e002f3c
0b06eabc
000760c3
601c0415
2ff3ff53
10f8501c
0000511c
8c0c740c
0080001c
44c62006
68c0301c
0016311c
b0c34664
64540007
8c0c740c
0080001c
44c62006
68c0301c
0016311c
c0c34664
740c06f2
0bc38c4c
09931cc3
20060bc3
0080201c
0891b0bc
20060cc3
0080201c
0891b0bc
253cadd7
1157fff0
141d6800
733c3350
8dc3528d
27d21dc3
68000dc3
3350141d
528d833c
278018c3
7e8021b7
23c33884
602761f7
901c2d35
911c10f8
19c30000
8c0c640c
329702c3
301c4066
311c68c0
46640016
4026a0c3
00074237
09c31d94
8c4c600c
1ac30bc3
301c44c6
311c68c0
46640016
640c19c3
0cc38c4c
44c61ac3
68c0301c
0016311c
d0664664
40062113
af3c4237
3ac30e70
62776e80
978493c3
1f5c0ac3
25c30921
0891b0bc
01538006
315704c3
0a7c6ebc
44222097
46212257
47e48025
8006f674
04c30153
6ebc1dc3
20d70a7c
19c34422
80254621
f67448e4
0e171513
31970037
12172077
41d71ac3
84bc3bc3
60c30b07
63dc0007
4006000a
6e170133
3230341d
21a20bc3
21210cc3
6dd74025
20e403c3
09c3f574
0ae25ebc
d24603d2
09c30293
4dd71cc3
0ae4e8bc
d22603d2
09c30193
29c32026
0aed86bc
b4dc0007
c3f2000a
0b7376c3
0cc00f3c
0ae27ebc
20060f33
20772037
18c30dc3
32c34006
0ae2a4bc
d24603d2
425709d3
0dc3ab80
4dd715c3
0ae4e8bc
0007d226
0dc33694
28c319c3
0ae67abc
d1a60177
2d940007
18bc08c3
40c30ae3
0007d1e6
4dd72674
0ef442e4
1f3c08c3
60bc02b0
60c30af2
1f3c05c3
4dd702c0
08cbb0bc
42e402d3
05c30f15
00a13f5c
4a2013c3
0891b0bc
7c000dd7
08c36e20
29804257
08c30073
60bc15c3
60c30af2
7ebc0dc3
08c30ae2
0ae27ebc
0774c007
fc000dd7
21c32197
a87472e4
2e1711d7
0b06d2bc
011740c3
24c31bc3
08cbb0bc
6e006117
11d76137
11f70220
7ebc09c3
00f30ae2
0cc09f3c
0bc0df3c
0ac08f3c
21c331d7
06dc4007
6217fff5
301c6fd2
311c10f8
6c0c0000
0ac38c4c
40663297
68c0301c
0016311c
501c4664
511c10f8
740c0000
0bc38c4c
44c62006
68c0301c
0016311c
740c4664
0cc38c4c
44c62006
68c0301c
0016311c
00734664
eb33d1a6
3a9606c3
0f56fc76
00000804
fa961016
80378217
80778257
80b78297
80f782d7
81378317
81778006
0b0836bc
08560696
00000804
3f36f016
fde0f21c
61c3a0c3
607782c3
12a49f5c
12c4bf5c
d8bc0bc3
c0c30b06
ff53501c
33dc0007
301c0008
311c10f8
6c0c0000
08068c0c
44c62006
68d4301c
0016311c
70c34664
0007b066
4f3c7054
04c30080
26c31bc3
26bc38c3
d0c30b1d
0001801c
0007b4c3
0a535054
20570bc3
12642f5c
0b1d14bc
000750c3
83064a94
408d283c
3f5c4037
3f5c0001
0bc310fd
21f01f3c
14bc4026
50c30b1d
39940007
9f079f05
0bc3ee94
04bc17c3
50c30b1d
2f940007
1cc309c3
0b06d2bc
0ac360c3
26c317c3
08cbb0bc
02d38026
17c30bc3
14bc2cc3
50c30b1d
1b940007
17c30bc3
0b1d04bc
000750c3
0ac31494
26c317c3
0b0696bc
3f5c8025
23c31284
e77442e4
96a4a684
0001821c
600739c3
5dc3b094
10f8301c
0000311c
8c4c6c0c
200607c3
301c44c6
311c68d4
46640016
f21c05c3
fc760220
08040f56
213cfe96
0080fff0
105c01f3
31c3fff9
60376025
00011f5c
3f5c2077
303c0021
24f2ffde
40075fe5
0296f115
00000804
0136f016
60c3fe96
23c342c3
2c542007
2a546007
281412e4
fff0513c
11002080
01b38006
87c3e409
8784e009
80374884
00017f5c
8017e40d
bfe58832
3fe55fe5
40071fe5
1a80f015
e0090193
80779380
00213f5c
ffdf303c
473ce057
bfe5820b
a00783d2
0296f315
0f568076
00000804
61c3f016
108c523c
701c8006
711c10fc
00d30000
6cac7c0c
1a613664
45e48085
0006fa14
08040f56
3f36f016
71c3d996
3f5c42c3
bf5c003d
af5c0684
323c06a4
6977180c
10bc03c3
09770b06
343c4006
62d201f4
343c4026
92c3288c
40269384
04dd2f5c
5f3cc006
df3c0080
cf3c0940
8f3c0070
0a330740
bebc05c3
00070b16
05c35594
09b01f3c
f6bc4026
00070b16
05c34d94
40861dc3
0b16f6bc
46940007
00393f5c
08546087
1cc305c3
f6bc4026
00070b16
05c33b94
4cd72c97
0b16f6bc
34940007
4ad22bc3
68d23ac3
1bc305c3
f6bc2ac3
00070b16
05c32994
3abc18c3
00070b17
84072394
07c30935
440618c3
08cbb0bc
e4059c05
07c300d3
24c318c3
08cbb0bc
2f5cc025
32c304d9
60376025
00011f5c
04dd1f5c
af7469e4
07400f3c
b8bc2406
00060b06
00460053
fc762796
08040f56
0136f016
70c3fa96
52c341c3
200663c3
b0bc4f06
873c0891
80370080
c0b7a077
60f76317
18c307c3
608646e6
0b0ae6bc
00070137
8f5c1a94
86e60007
00b78077
07c300f7
03f0173c
4f5c24c3
34c30081
0b0ae6bc
09f20177
7c0f6026
3f5c1c2f
375c00a1
005303b5
06960046
0f568076
00000804
ec967016
503c40c3
6f3c0080
a0370190
607766e6
40f720b7
23c316c3
e6bc6026
01370b0a
23940007
16c305c3
b0bc46e6
06c308cb
b8bc26e6
a0370b06
a077a6e6
60b76117
04c360f7
03f0143c
5f5c25c3
35c30081
0b0ae6bc
09f20177
700f6026
3f5c102f
345c00a1
005303b5
14960046
08040e56
1f36f016
60c3ce96
52c371c3
42f213c3
4006a026
01f4353c
402662d2
288c353c
a384a2c3
06d04f3c
46e604c3
08cbb0bc
0000801c
4f3cb4c3
cf3c0a40
09130c40
bebc0fc3
00070b16
0fc34c94
46e61bc3
0b16f6bc
45940007
14c30fc3
0b173abc
3f940007
14c30cc3
b0bc4086
780c08cb
10356027
582c6c57
30e402c3
365c0b94
602703b1
00860394
402605b3
03b5265c
600600d3
03b5365c
182f0c57
1654e007
0d35a3e7
14c307c3
b0bc4406
bc0508cb
0bc3e405
82bc26e6
01130b0a
07c3a7d2
25c314c3
08cbb0bc
821ca006
8ae40001
0f3cb874
26e606d0
0b06b8bc
00530006
32960046
0f56f876
00000804
0136f016
60c3db96
e066600c
4240401c
000f411c
35e454c3
80664854
049d4f5c
503c68f7
35c30080
0b0be0bc
000770c3
0fc33c94
0b16bebc
33940007
1f3c0fc3
40260930
0b16f6bc
2b940007
15c30fc3
f6bc46e6
00070b16
8f3c2494
0fc306c0
3abc18c3
00070b17
05c31c94
28c326e6
9abc6406
05c30b0a
263c26e6
31c303f0
0b0a9abc
10bc08d7
3f3c0b06
033c0940
05c3fc7e
23c326e6
9abc6086
00530b0a
780ce046
780f6025
06c00f3c
b8bc2406
07c30b06
80762596
08040f56
40c31016
b8bc2f06
60060b06
51a203c3
602502a3
fc946f07
004602d2
08040856
0f36f016
71c3ff96
a3c382c3
0164bf5c
e2dc2007
2bc3000b
a2dc4007
303c000b
33c40b0d
f88c933c
65d239c3
40072ac3
000af2dc
331c6317
d4dc0080
301c000a
311c10f8
6c0c0000
0f068c0c
44062006
6c30301c
0016311c
60c34664
0007b066
0009b2dc
60376006
28c317c3
0b0b6cbc
79940007
101c07c3
111c68e0
46060016
08cbeabc
17940007
6960001c
0016011c
0080163c
eabc46e6
000708cb
001c7c94
011c6998
163c0016
46e603f0
08cbeabc
71940007
101c07c3
111c6910
46060016
08cbeabc
17940007
69d0001c
0016011c
0080163c
eabc46e6
000708cb
001c5c94
011c6a08
163c0016
46e603f0
08cbeabc
51940007
48d229c3
1ac306c3
a6bc4297
00070b0b
07c33094
6940101c
0016111c
eabc4406
000708cb
001c1794
011c6a40
163c0016
46e60080
08cbeabc
33940007
6a78001c
0016011c
03f0163c
eabc46e6
000708cb
06c32894
201c1bc3
56bc0080
09f20b0c
1bc306c3
0080201c
0b0c56bc
02d250c3
06c3bfe6
0b0cb4bc
bfe602d2
10f8301c
0000311c
8c4c6c0c
200606c3
301c4406
311c6c30
46640016
501c00b3
0053ff53
05c3bfe6
f0760196
08040f56
60c37016
ff53501c
1e540007
501c000c
0007ff53
b4bc1754
50c30b0c
501c03d2
301cff39
311c10f8
6c0c0000
180c8c4c
4406384c
6c44301c
0016311c
60064664
6006780f
05c3798d
08040e56
fd96f016
301c60c3
311c10f8
6c0c0000
001c8c0c
20060080
301c44c6
311c6c50
46640016
b06670c3
47540007
1c54c007
60376406
301c0077
60b70080
101c0026
111c6ab0
46060016
6ae0301c
0016311c
0b0cc4bc
000750c3
07c32294
6b00101c
0016111c
c03702d3
301c0077
60b70080
101c06c3
111c6b80
46060016
c4bc36c3
50c30b0c
07c30cf2
6bb0101c
0016111c
0080201c
0b06c0bc
bfe602d2
10f8301c
0000311c
8c4c6c0c
200607c3
301c44c6
311c6c50
46640016
039605c3
08040f56
0136f016
50c3f896
82c371c3
51540007
4f542007
011c0006
30c30001
49b423e4
401cd589
c027ff39
140c4694
0b0c56bc
006740c3
06c33194
0b0dbabc
2f940007
10fc301c
0000311c
6d0c6c0c
80463664
31940007
0040053c
44061fc3
0b0ad2bc
15940007
1fc3140c
a6bc4406
10c30b0b
140c0ef2
56bc21c3
40c30b0c
140c09f2
28c317c3
0b0c56bc
005340c3
0fc38046
b8bc2406
8fd20b06
06948087
758d6066
ff2f401c
00460113
401c158d
0073ff39
ff53401c
089604c3
0f568076
00000804
1abc4026
08040b0e
f2967016
301c50c3
6077ff53
58540007
0006204f
0b0dbabc
3f940007
10f8301c
0000311c
8c0c6c0c
344c0f06
301c4406
311c6c68
46640016
5066140f
00074077
6f3c1e54
053c0080
16c30040
d2bc4606
40c30b0a
11940007
0037740c
16c303c3
34c34606
0b0b6cbc
07f210c3
21c3140c
0b0c56bc
00730077
60776046
00800f3c
b8bc2606
40570b06
602644f2
0313758d
32c34057
07946087
558d4066
ff2f201c
01d34077
23c36057
08944047
00213f5c
301c758d
6077ff39
40460073
0057558d
0e560e96
00000804
7ebc2006
08040b0e
ff53301c
18540007
305c7fe6
60060407
0447305c
0427105c
0467305c
0487305c
04a5305c
60ef6006
61ef606f
62ef616f
636f626f
03c363ef
00000804
e6bc5fc6
08040b0e
0736f016
73c3a2c3
813c7264
2147ff60
801c03b4
3ac30000
24f262d2
ff53001c
905c0633
60c30001
fff0413c
009e563c
202620c3
0b9471e4
14e417c3
60490e34
00252025
00ff331c
00f3f954
053414e4
20256849
7bf24025
055414e4
235c7880
4ef2fff9
570310a0
39c425c4
7f3232a3
06b408e4
788065f2
680f2ac3
001c0073
e076ff37
08040f56
0ae318bc
00000804
0736f016
81c360c3
a3c352c3
01049f5c
2c540007
2a542007
28544007
26546007
200719c3
403c2354
04c30100
0ae318bc
540c70c3
03e432c3
04c31cb4
60bc18c3
00070af2
f40f1894
4cbc06c3
40c30b0f
440c19c3
03e432c3
06c30cb4
60bc1ac3
09f20af2
840f19c3
001c00d3
0073ff53
ff7d001c
0f56e076
00000804
0336f016
90c3ff96
52c341c3
01011f5c
00072037
80074454
40074254
60074054
40063e54
75c3540d
fff0633c
00013f5c
00de373c
0e942027
0020343c
321463e4
073c7a20
3fe60010
ffe0233c
0891b0bc
343c0353
63e40010
34e32514
868483c3
173c0257
28c30010
0b0e1abc
602625c3
035308d2
23f22849
284d2026
40256025
f91438e4
7d807a20
235c4006
03c3fffd
24c319c3
08cbb0bc
00d30006
ff53001c
001c0073
0196ff37
0f56c076
00000804
3f36f016
01f7e696
a2c321b7
f0bc6177
70c30b23
63dc0007
9a3c0009
931c0040
08b40044
02406f3c
801c8006
08e40044
87c31835
023479e4
301c89c3
311c10f8
6c0c0000
08c38c0c
44c62997
6c84301c
0016311c
60c34664
03f28026
0e53f066
22372006
2ac3b1c3
133c7900
20770010
0020d33c
0030c33c
219706c3
b0bc2ac3
421708cb
41375832
00815f5c
b9a13ac3
30322217
3f5c20f7
40570061
a217680d
a0b7a832
00412f5c
440d1dc3
01015f5c
ac0d3cc3
00078f5c
16c301d7
36c329c3
0b257cbc
05f250c3
21573bc3
03134580
800770c3
301c3754
311c10f8
6c0c0000
06c38c4c
44c62997
6c84301c
0016311c
75c34664
b82204f3
6025a821
07e40025
a9570515
31e415c3
4957f714
35e452c3
22170734
402521c3
b3c34237
74c3f5d3
10548007
10f8301c
0000311c
8c4c6c0c
299706c3
301c44c6
311c6c84
46640016
07c3e006
fc761a96
08040f56
fe967016
a1d78197
15540047
04d40047
06940027
00670193
03471254
001c0454
0253ff53
a0778037
01930086
a0778037
011300a6
a0778037
009300c6
a0778037
e6bc00e6
02960b0f
08040e56
3f36f016
0177f896
c2c391c3
e5d76137
0304af5c
0324bf5c
601ce7f2
0ac3ff7c
64dc0007
0557001a
0b23f0bc
000760c3
0019f3dc
10f8501c
0000511c
8c0c740c
44c61bc3
6c78301c
0016311c
80c34664
17540007
8c0c740c
1bc306c3
301c44c6
311c6c78
46640016
0df2d0c3
8c4c740c
1bc308c3
301c44c6
311c6c78
46640016
2ed3d066
0557c037
2ac317c3
7cbc38c3
70c30b25
740c0dd2
08c38c4c
44c61bc3
6c78301c
0016311c
740c4664
363c1b73
61b70010
81176112
30e404c3
163c09b4
41170b0c
7fc532c3
93e46c80
740c1835
08c38c4c
44c61bc3
6c78301c
0016311c
740c4664
0dc38c4c
44c61bc3
6c78301c
0016311c
601c4664
2753ff53
20c30117
183429e4
8c4c740c
1bc308c3
301c44c6
311c6c78
46640016
8c4c740c
1bc30dc3
301c44c6
311c6c78
46640016
ff7c601c
811723f3
39a434c3
fff0533c
ffe0233c
0cc3e880
04c38180
29c32157
08cbb0bc
1cc34026
353c46a1
00d3fff0
045c0006
7fe5fffd
9fe5ffe5
02f4e007
6f2078f2
2cc36025
18c30980
b0bc26c3
051708cb
26c31dc3
0b0e1abc
901c01f7
911c10f8
00070000
49c31954
8c4c700c
1bc308c3
301c44c6
311c6c78
46640016
600c09c3
0dc38c4c
44c61bc3
6c78301c
0016311c
c1d74664
21171ab3
7fe531c3
a6a4a3c3
700c49c3
0ac38c0c
41461bc3
6c78301c
0016311c
50c34664
11940007
600c09c3
08c38c4c
44c61bc3
6c78301c
0016311c
19c34664
8c4c640c
e6930dc3
00e12f5c
2ac312c3
0891b0bc
0007af5c
0027bf5c
1dc30597
35c326c3
0b108cbc
000770c3
49c32454
8c4c700c
1bc305c3
301c4146
311c6c78
46640016
600c09c3
08c38c4c
44c61bc3
6c78301c
0016311c
19c34664
8c4c640c
1bc30dc3
301c44c6
311c6c78
46640016
0f9367c3
6b002cc3
01734197
14c38c09
14039422
1f5c20f7
2c0d0061
40250025
14c38117
043421e4
0ae46025
701cf014
711c10f8
7c0c0000
05c38c4c
41461bc3
6c78301c
0016311c
20064664
200d0cc3
0010363c
bf5cc037
05970027
29802cc3
3c3c2ac3
8cbc0010
50c30b10
602620c3
25540007
8c4c7c0c
1bc308c3
301c44c6
311c6c78
46640016
8c4c7c0c
1bc30dc3
301c44c6
311c6c78
46640016
05d365c3
11224dc3
4cc310c3
40c311a2
20b71403
00411f5c
21a10cc3
60254025
04c38197
033430e4
ed7426e4
10f8501c
0000511c
8c4c740c
1bc308c3
301c44c6
311c6c78
46640016
8c4c740c
1bc30dc3
301c44c6
311c6c78
46640016
06c3c006
fc760896
08040f56
f896f016
a3d7c397
01a14f5c
a6d281f7
ff37401c
1c94a027
4f5c0133
4f5c00e1
c0770005
0b0f8ebc
7f5c0253
7f5c00e1
c0770005
80b78417
e0f7e457
81378497
e177e4d7
81b78517
0b10b2bc
04c340c3
0f560896
00000804
3f36f016
80c3ea96
4177a1c3
bf5c6137
28970484
501c27f2
48d7ff7c
a4dc4007
0117000b
0b23f0bc
000770c3
000b13dc
0010903c
080c393c
a0dca3e4
c01c000a
c11c10f8
1cc30000
8c0c640c
1bc30ac3
301c44c6
311c6ca0
46640016
b06660c3
82dc0007
20060009
b0bc2ac3
d8c30891
3a3cd984
93c3fff0
e03797a4
0027bf5c
1dc30857
36c329c3
0b108cbc
03f250c3
021336c3
640c1cc3
002504b3
882228c3
8c0914c3
120324c3
4f5c20f7
433c0061
07e400df
9b80f314
00079f5c
0027bf5c
16c30857
34c327c3
0b108cbc
05f250c3
4f8038c3
033334c3
10f8301c
0000311c
8c4c6c0c
200606c3
301c44c6
311c6ca0
46640016
8c2209f3
880914c3
20b71403
00411f5c
0025280d
09e44025
301cf514
311c10f8
6c0c0000
06c38c4c
44c61bc3
6ca0301c
0016311c
373c4664
433c080c
18c30010
00534580
4ae48025
323c0434
7bd2009e
01806f3c
0117e037
48d72897
7cbc36c3
50c30b25
1c940007
16c30dc3
c0bc27c3
18c30b06
32c34622
0001361c
6c802409
501c6c00
6cf2ff3f
0010243c
710048c3
640f2157
ad203ac3
501c0073
05c3ff53
fc761696
08040f56
fb963016
32648217
86d26137
ff37301c
14948027
4f5c00f3
34c30081
0b0f08bc
a2970193
62d7a037
83176077
a35780b7
6257a0f7
0b129abc
03c330c3
0c560596
00000804
50c33016
2a540007
0464005c
26540007
04a1255c
1d544007
0404355c
60277fc5
155c05b4
b8bc0484
301c0b06
311c10f8
6c0c0000
055c8c4c
155c0464
41460424
6cb0301c
0016311c
60064664
04a5355c
255c4006
255c0467
0c560487
00000804
0f36f016
80c3f496
a2c391c3
a557b3c3
7f3cc597
07c30200
0ae25ebc
00079246
0009b4dc
18c307c3
e8bc29c3
92260ae4
e4dc0007
a0070008
a0270574
a0675cf4
401c04f4
1093ff7e
01005f3c
5ebc05c3
92460ae2
7c940007
5ebc0fc3
06d20ae2
7ebc05c3
92460ae2
963c0e73
07c30300
0500163c
35c329c3
0afbd4bc
30940007
0400863c
163c07c3
28c30600
d4bc3fc3
00070afb
05c32594
27c31fc3
0ae698bc
000791c6
5f3c1e94
05c30200
0700163c
35c329c3
0af574bc
00079166
05c31294
25c318c3
0aefaabc
0bf29186
1fc305c3
7abc25c3
40c30ae6
91a604d2
92060053
01000f3c
0ae27ebc
7ebc0fc3
80070ae2
01732f94
163c07c3
26c30100
d4bc37c3
92060afb
24940007
4cbc06c3
50c30b0f
ff7d401c
440c1bc3
03e432c3
0f3c19b4
18bc0200
01130ae3
1ac34006
0001a21c
00df213c
05e40025
1bc3f814
0f3ca40f
1ac30200
0af260bc
02d240c3
0f3c91e6
7ebc0200
04c30ae2
f0760c96
08040f56
0336f016
8f5cfd96
a2d70144
1454a007
12540007
10542007
6ed24fd2
8cd28c0c
ffff831c
8f5c0954
a0770007
a0b7a317
0b13babc
001c0073
0396ff53
0f56c076
00000804
0736f016
80c3f796
72c361c3
a45793c3
0324af5c
02612f5c
00074237
20075e54
e0075c54
a0075a54
05c35854
0b0f4cbc
09e440c3
001c55d4
8147ff16
343c53f4
63e4ff50
355c4db4
60470444
60472954
600704d4
00730715
34546067
ff40001c
60460713
0447355c
01012f5c
00052f5c
0027af5c
60b76517
40f74557
61376597
417745d7
61b76617
0424255c
08c341f7
27c316c3
6ebc34c3
00070b12
40661874
0447255c
933c35c3
4497487e
a0774037
0047af5c
14c307c3
6abc27c3
00070b14
40060674
0447255c
0484055c
0a541287
255c4006
00d30447
ff53001c
001c0073
0996ff7d
0f56e076
00000804
f7961016
803782d7
80778046
4f5c8026
80060045
813780f7
81b78177
831781f7
8cbc8237
09960b14
08040856
f7961016
803782d7
80778006
4f5c8046
83570045
839780f7
83d78137
84178177
845781b7
831781f7
8cbc8237
09960b14
08040856
f7963016
80378317
80778006
5f5ca046
80f70045
81778137
81f781b7
82378357
0b148cbc
0c560996
00000804
0736f016
80c3f896
72c361c3
9f5ca3c3
a4570204
02610f5c
28c301b7
92dc4007
20070009
000962dc
32dce007
a0070009
000902dc
0444355c
0c546087
03d46087
0fd369d2
415460a7
ff53401c
789460c7
40a60e33
0447255c
0464355c
70946007
0487655c
600739c3
301c1d94
311c10f8
6c0c0000
06c38c0c
0424155c
301c4146
311c6c8c
46640016
0467055c
455c8026
906604a5
56540007
26c318c3
08cbb0bc
755c0073
355c0467
04970464
a0770037
40b74657
16c303c3
353c23c3
6abc0900
40c30b14
39740007
02003f3c
433c8006
00c6fe7e
0447055c
0464255c
0484155c
80378517
00770557
80b78597
00f705d7
81378617
0424055c
02c30177
4f5c23c3
34c300c1
0b1368bc
800740c3
4ae410f4
21d70ed4
20542007
66f239c3
24c307c3
08cbb0bc
09c300f3
0093200f
14158007
60060093
0447355c
04949287
401c0213
4006ff40
0447255c
8abc05c3
00f30b13
ff53401c
401c0093
fdf3ff7d
089604c3
0f56e076
00000804
f6963016
80378006
a077a357
a0b7a026
00655f5c
81778137
81f781b7
82778237
0b1548bc
0c560a96
00000804
4037f696
60266077
3f5c60b7
60060065
61776137
61f761b7
62776237
31c320c3
0b1548bc
08040a96
f6963016
80378006
a077a357
a0b7a066
5f5ca046
a3970065
a3d7a137
a417a177
a457a1b7
a497a1f7
8277a237
0b1548bc
0c560a96
00000804
f6963016
80378006
a077a357
a0b7a066
5f5ca046
81370065
81b78177
823781f7
48bc8277
0a960b15
08040c56
4037f696
60666077
604660b7
00653f5c
613762d7
61776317
61b76357
61f76397
623763d7
62776006
31c320c3
0b1548bc
08040a96
4037f696
60666077
604660b7
00653f5c
61376006
61b76177
623761f7
20c36277
48bc31c3
0a960b15
00000804
40c31016
ff53301c
27540007
0b138abc
0404345c
19946027
0700043c
0afd36bc
0600043c
0afd36bc
0500043c
0afd36bc
0400043c
0afd36bc
0300043c
0afd36bc
0200043c
0afd36bc
0100043c
0ae27ebc
7ebc04c3
60060ae2
085603c3
00000804
01c330c3
023513e4
080403c3
e667201c
6a09211c
201c406f
211cae85
408fbb67
f372201c
3c6e211c
201c40af
211cf53a
40cfa54f
527f201c
510e211c
201c40ef
211c688c
410f9b05
d9ab201c
1f83211c
201c412f
211ccd19
414f5be0
400f4006
404f402f
080402c3
6500402c
32e4602f
604c0434
604f6025
00000804
3f36f016
50c3ff96
82c391c3
02c0a03c
00c0b03c
10f8d01c
0000d11c
10fcc01c
0000c11c
940c0533
480608c3
b8bc2a20
70c30b16
0e003ac3
27c319c3
08cbb0bc
dc80340c
c807d40f
1dc31594
1cc3640c
28a9440c
00051f5c
0ac38d6c
40461bc3
46646006
0cf240c3
16c305c3
0b16ecbc
9784940f
28c387a4
d6944007
04c348c3
fc760196
08040f56
0136f016
50c3ff96
703c81c3
200c02c0
0b16ecbc
1006740c
60251da1
6707740f
88062035
20061d80
b0bc51a0
25c30891
067f423c
10f8301c
0000311c
301c2c0c
311c10fc
6c0c0000
0f5c0ca9
856c0005
12c307c3
60064046
00074664
140f4c94
1d00540c
67062006
b0bc4d20
744c0891
180c133c
323c542c
6580e88c
323c744f
742f180c
0380073c
0080153c
b0bc4086
073c08cb
153c03c0
40860040
08cbb0bc
0640353c
13c303c3
24bc4106
653c0b06
301c00c0
311c10f8
4c0c0000
10fc301c
0000311c
2ca96c0c
00051f5c
07c3896c
404616c3
46646006
06c30ef2
440616c3
0b0624bc
16c308c3
b0bc4406
05c308cb
0b16bebc
80760196
08040f56
01c330c3
023513e4
080403c3
c908201c
f3bc211c
201c406f
211ce667
408f6a09
a73b201c
84ca211c
201c40af
211cae85
40cfbb67
f82b201c
fe94211c
201c40ef
211cf372
410f3c6e
36f1201c
5f1d211c
201c412f
211cf53a
414fa54f
82d1201c
ade6211c
201c416f
211c527f
418f510e
6c1f201c
2b3e211c
201c41af
211c688c
41cf9b05
bd6b201c
fb41211c
201c41ef
211cd9ab
420f1f83
2179201c
137e211c
201c422f
211ccd19
424f5be0
400f4006
404f402f
080402c3
6500402c
32e4602f
604c0434
604f6025
00000804
9ed8201c
c105211c
201c406f
211c9d5d
408fcbbb
d507201c
367c211c
201c40af
211c292a
40cf629a
dd17201c
3070211c
201c40ef
211c015a
410f9159
5939201c
f70e211c
201c412f
211cecd8
414f152f
0b31201c
ffc0211c
201c416f
211c2667
418f6733
1511201c
6858211c
201c41af
211c4a87
41cf8eb4
8fa7201c
64f9211c
201c41ef
211c2e0d
420fdb0c
4fa4201c
befa211c
201c422f
211c481d
424f47b5
400f4006
404f402f
080402c3
6500402c
32e4602f
604c0434
604f6025
00000804
0136f016
50c3ff96
703c81c3
200c04c0
0b1874bc
1006740c
60251da1
6e07740f
401c2135
1d800080
51a02006
0891b0bc
423c25c3
301c067f
311c10f8
2c0c0000
10fc301c
0000311c
0ca96c0c
00050f5c
07c3856c
406612c3
46646006
46940007
540c140f
20061d00
4d206e06
0891b0bc
133c744c
542c180c
e88c323c
744f6580
542f4312
05e7355c
155c2006
255c0607
155c0627
353c0647
03c30bc0
420613c3
0b0672bc
10f8301c
0000311c
653c4c0c
301c00c0
311c10fc
6c0c0000
0f5c0ca9
896c0005
16c307c3
60064066
0ef24664
16c306c3
72bc4606
08c30b06
460616c3
08cbb0bc
1ebc05c3
01960b18
0f568076
00000804
3f36f016
50c3ff96
82c391c3
04c0a03c
00c0b03c
10f8d01c
0000d11c
10fcc01c
0000c11c
940c0573
201c08c3
2a200080
0b17b8bc
3ac370c3
19c30e00
b0bc27c3
340c08cb
d40fdc80
0080631c
1dc31594
1cc3640c
28a9440c
00051f5c
0ac38d6c
40661bc3
46646006
0cf240c3
16c305c3
0b1874bc
9784940f
28c387a4
d4944007
04c348c3
fc760196
08040f56
0136f016
50c3ff96
703c81c3
200c04c0
0b1814bc
1006740c
60251da1
6e07740f
401c2135
1d800080
51a02006
0891b0bc
423c25c3
301c067f
311c10f8
2c0c0000
10fc301c
0000311c
0ca96c0c
00050f5c
07c3856c
408612c3
46646006
46940007
540c140f
20061d00
4d206e06
0891b0bc
133c744c
542c180c
e88c323c
744f6580
542f4312
05e7355c
155c2006
255c0607
155c0627
353c0647
03c30bc0
420613c3
0b0672bc
10f8301c
0000311c
653c4c0c
301c00c0
311c10fc
6c0c0000
0f5c0ca9
896c0005
16c307c3
60064086
0ef24664
16c306c3
72bc4806
08c30b06
480616c3
08cbb0bc
bebc05c3
01960b17
0f568076
00000804
3f36f016
50c3ff96
82c391c3
04c0a03c
00c0b03c
10f8d01c
0000d11c
10fcc01c
0000c11c
940c0573
201c08c3
2a200080
0b17b8bc
3ac370c3
19c30e00
b0bc27c3
340c08cb
d40fdc80
0080631c
1dc31594
1cc3640c
28a9440c
00051f5c
0ac38d6c
40861bc3
46646006
0cf240c3
16c305c3
0b1814bc
9784940f
28c387a4
d4944007
04c348c3
fc760196
08040f56
01c330c3
023513e4
080403c3
2301201c
6745211c
201c426f
211cab89
428fefcd
dcfe201c
98ba211c
201c42af
211c5476
42cf1032
e1f0201c
c3d2211c
400642ef
402f400f
02c3404f
00000804
6500402c
32e4602f
604c0434
604f6025
00000804
1f36f016
50c3ff96
72c381c3
00c0903c
04c0a03c
0040c01c
10fcb01c
0000b11c
940c04d3
2cc307c3
febc2a20
60c30b19
0e0039c3
26c318c3
08cbb0bc
9900540c
8807940f
2bc31294
4ca9680c
00052f5c
1ac309c3
32c34006
087d86bc
14c305c3
0b1a24bc
740f6006
ff208684
da94e007
019607c3
0f56f876
00000804
ff96f016
71c350c3
00c0603c
24bc200c
740c0b1a
39a13006
740f6025
1a356707
19808806
51a02006
0891b0bc
423c25c3
301c267f
311c10fc
6c0c0000
1f5c2ca9
06c30005
400612c3
86bc32c3
4006087d
540c540f
20061900
4d206706
0891b0bc
133c744c
542c180c
e88c323c
744f6580
180c323c
063c742f
153c0380
40860080
08cbb0bc
03c0063c
0040153c
b0bc4086
353c08cb
03c30440
410613c3
0b0624bc
04c0453c
10fc301c
0000311c
2ca96c0c
00051f5c
14c306c3
32c34006
087d86bc
14c304c3
24bc4286
07c30b06
428614c3
08cbb0bc
04bc05c3
01960b1a
08040f56
13cc301c
0000311c
00060c0f
00000804
401c1016
411c10fc
700c0000
36646ccc
602730c3
700c1754
20072c89
6c0c3754
0bc1035c
035c10c3
203c0bc9
135c40ac
213c0bd1
035c812c
303c0bd9
6027c12c
301c2594
311c13d0
6c0c0000
1e546047
14946027
13cc301c
0000311c
80078c0c
00061754
13d8301c
0000311c
201c2c0c
211c13dc
46640000
6af20173
13d4301c
0000311c
60276c0c
00060394
1fe60053
08040856
301c1016
311c13d0
40060000
301c4c0f
311c13d4
40260000
301c4c0f
311c10f8
6c0c0000
001c6c8c
011c13dc
36640000
13d8401c
0000411c
0cf2100f
10fc301c
0000311c
4c896c0c
6cec4bd2
100f3664
301c07d2
311c13d0
40260000
301c00d3
311c13d0
40460000
301c4c0f
311c13d4
40060000
08564c0f
00000804
0b1b2ebc
00000804
0136f016
61c350c3
83c372c3
0b1ae4bc
ff3b301c
301c0df2
311c10fc
6c0c0000
05c38f0c
27c316c3
466438c3
03c330c3
0f568076
00000804
40c33016
e4bc51c3
301c0b1a
0bf2ff3b
10fc301c
0000311c
6f2c6c0c
15c304c3
30c33664
0c5603c3
00000804
0136f016
61c350c3
83c372c3
0b1ae4bc
ff3b301c
301c0df2
311c10fc
6c0c0000
05c38f6c
27c316c3
466438c3
03c330c3
0f568076
00000804
0136f016
61c350c3
83c372c3
0b1ae4bc
ff3b301c
301c0df2
311c10fc
6c0c0000
05c38f4c
27c316c3
466438c3
03c330c3
0f568076
00000804
fd96f016
51c340c3
73c362c3
0b1ae4bc
ff3b301c
62170ef2
62576037
62976077
04c360b7
26c315c3
c4bc37c3
30c30b0c
039603c3
08040f56
40c37016
62c351c3
0b1ae4bc
ff3b301c
04c307f2
26c315c3
0b0e1abc
03c330c3
08040e56
40c31016
0b1ae4bc
ff3b301c
04c305f2
0b0d94bc
03c330c3
08040856
40c31016
0b1ae4bc
ff3b301c
04c305f2
0b0ee2bc
03c330c3
08040856
40c3f016
62c351c3
e4bc73c3
301c0b1a
08f2ff3b
15c304c3
37c326c3
0ac042bc
03c330c3
08040f56
40c3f016
62c351c3
e4bc73c3
301c0b1a
08f2ff3b
15c304c3
37c326c3
0abeb4bc
03c330c3
08040f56
40c31016
0b1ae4bc
ff3b301c
04c305f2
0b0f4cbc
03c330c3
08040856
ff96f016
51c340c3
73c362c3
0b1ae4bc
ff3b301c
61970af2
04c36037
26c315c3
fcbc37c3
30c30b15
019603c3
08040f56
40c3f016
62c351c3
e4bc73c3
301c0b1a
08f2ff3b
15c304c3
37c326c3
0b1612bc
03c330c3
08040f56
fe96f016
51c340c3
73c362c3
0b1ae4bc
ff3b301c
61d70cf2
62176037
04c36077
26c315c3
02bc37c3
30c30b15
029603c3
08040f56
ff96f016
51c340c3
73c362c3
0b1ae4bc
ff3b301c
61970af2
04c36037
26c315c3
42bc37c3
30c30b16
019603c3
08040f56
40c3f016
62c351c3
e4bc73c3
301c0b1a
08f2ff3b
15c304c3
37c326c3
0b1672bc
03c330c3
08040f56
fe96f016
51c340c3
73c362c3
0b1ae4bc
ff3b301c
61d70cf2
62176037
04c36077
26c315c3
32bc37c3
30c30b15
029603c3
08040f56
40c31016
0b1ae4bc
ff3b301c
04c305f2
0b1688bc
03c330c3
08040856
40c33016
e4bc51c3
301c0b1a
06f2ff3b
15c304c3
0b0f04bc
03c330c3
08040c56
40c33016
e4bc51c3
301c0b1a
06f2ff3b
15c304c3
0adf9abc
03c330c3
08040c56
40c37016
62c351c3
0b1ae4bc
ff3b301c
04c307f2
26c315c3
0ae042bc
03c330c3
08040e56
40c3f016
62c351c3
e4bc73c3
301c0b1a
08f2ff3b
15c304c3
37c326c3
0ae0bcbc
03c330c3
08040f56
40c33016
e4bc51c3
301c0b1a
06f2ff3b
15c304c3
0b187ebc
03c330c3
08040c56
40c37016
62c351c3
0b1ae4bc
ff3b301c
04c307f2
26c315c3
0b18f8bc
03c330c3
08040e56
40c31016
0b1ae4bc
ff3b301c
04c305f2
0b181ebc
03c330c3
08040856
40c33016
e4bc51c3
301c0b1a
06f2ff3b
15c304c3
0b193ebc
03c330c3
08040c56
40c37016
62c351c3
0b1ae4bc
ff3b301c
04c307f2
26c315c3
0b19b8bc
03c330c3
08040e56
40c31016
0b1ae4bc
ff3b301c
04c305f2
0b17bebc
03c330c3
08040856
40c33016
e4bc51c3
301c0b1a
06f2ff3b
15c304c3
0b173abc
03c330c3
08040c56
40c37016
62c351c3
0b1ae4bc
ff3b301c
04c307f2
26c315c3
0b16f6bc
03c330c3
08040e56
40c31016
0b1ae4bc
ff3b301c
04c305f2
0b16bebc
03c330c3
08040856
40c33016
e4bc51c3
301c0b1a
06f2ff3b
15c304c3
0b1a6cbc
03c330c3
08040c56
40c37016
62c351c3
0b1ae4bc
ff3b301c
04c307f2
26c315c3
0b1a2ebc
03c330c3
08040e56
40c31016
0b1ae4bc
ff3b301c
04c305f2
0b1a04bc
03c330c3
08040856
fa96f016
51c340c3
73c362c3
0b1ae4bc
ff3b301c
14940007
603762d7
60776317
60b76357
60f76397
613763d7
61776417
15c304c3
37c326c3
0a9f5cbc
03c330c3
0f560696
00000804
fa96f016
51c340c3
73c362c3
0b1ae4bc
ff3b301c
14940007
603762d7
60776317
60b76357
60f76397
613763d7
61776417
15c304c3
37c326c3
0a9ff6bc
03c330c3
0f560696
00000804
40c37016
62c351c3
0b1ae4bc
ff3b301c
04c307f2
26c315c3
0aa098bc
03c330c3
08040e56
40c3f016
62c351c3
e4bc73c3
301c0b1a
08f2ff3b
15c304c3
37c326c3
0a9b58bc
03c330c3
08040f56
40c3f016
62c351c3
e4bc73c3
301c0b1a
08f2ff3b
15c304c3
37c326c3
0a9ba8bc
03c330c3
08040f56
40c33016
e4bc51c3
301c0b1a
06f2ff3b
15c304c3
0a9a2abc
03c330c3
08040c56
ff96f016
51c340c3
73c362c3
0b1ae4bc
ff3b301c
61970af2
04c36037
26c315c3
f6bc37c3
30c30a99
019603c3
08040f56
0336f016
82c371c3
501c93c3
511c10f8
740c0000
7ca4601c
0016611c
20068c4c
36c344c6
740c4664
07c38c4c
44c62006
466436c3
8c4c740c
200608c3
36c344c6
740c4664
09c38c4c
44c62006
466436c3
8c4c740c
200601d7
36c344c6
c0764664
08040f56
3f36f016
b0c38996
d2c3c1c3
6f5c6077
af5c1063
301c10a3
311c10f8
6c0c0000
001c8c0c
20060098
301c44c6
311c7794
46640016
506650c3
6a540007
19c07f3c
280607c3
08cb9cbc
13809f3c
2c8609c3
08cb9cbc
0d408f3c
2c8608c3
08cb9cbc
101c05c3
9cbc0098
4f3c08cb
04c30080
00cc101c
08cb9cbc
200605c3
0b1cf4bc
ff47201c
44940007
0f5ca037
16c31044
10842f5c
2ebc3ac3
60c30abe
05c307d2
0b1ce6bc
ff47201c
04c30673
0b1d8cbc
1bc304c3
7abc2cc3
04c30b1d
6abc17c3
00860b1d
0aa532bc
09c330c3
480617c3
0ab594bc
a03740c3
20570dc3
6c8628c3
0b1c5abc
05c370c3
0b1ce6bc
05c3c037
26c316c3
a4bc36c3
74e40b1e
08c30894
27c319c3
08cbeabc
02d220c3
02c35fe6
fc767796
08040f56
3f36f016
60c3ff96
82c371c3
af5c93c3
bf5c0184
cf5c01a4
df5c01c4
313c01e4
33c40b0d
f88c533c
33540007
3154a007
2f544007
08920ebc
784b203c
4c0f38c3
10f8301c
0000311c
8c0c6c0c
200602c3
301c44c6
311c7c94
46640016
90661c0f
f2dc0007
06c3000f
08920ebc
336430c3
13c306c3
38c35c0c
0ac9dabc
09d240c3
a0067c0c
03c3a037
25c315c3
1cb335c3
0b0d3a3c
633c33c4
29c3f88c
3e544007
3c54c007
60073bc3
09c33954
08920ebc
784b203c
4c0f3bc3
10f8301c
0000311c
8c0c6c0c
200602c3
301c44c6
311c7c94
46640016
080f2ac3
05c309f2
1c0ca2d2
60376006
23c313c3
09c312d3
08920ebc
336430c3
13c309c3
4c0c3ac3
dabc3bc3
40c30ac9
05c30bd2
1c0ca2d2
740c5ac3
40374006
32c313c3
3d3c1413
33c40b0d
f88c833c
60073cc3
28c34754
44544007
60076417
0cc34154
08920ebc
784b203c
4c0f6417
10f8301c
0000311c
8c0c6c0c
200602c3
301c44c6
311c7c94
46640016
080f2dc3
05c30df2
1c0ca2d2
c3d216c3
2c0c3ac3
a037a006
35c325c3
0cc30993
08920ebc
336430c3
13c30cc3
4c0c3dc3
dabc6417
40c30ac9
05c30fd2
1c0ca2d2
c3d216c3
340c5ac3
680c2dc3
a037a006
35c323c3
44570a53
52544007
60076497
44d74f54
4c544007
0ebc0457
203c0892
64d7784b
301c4c0f
311c10f8
6c0c0000
02c38c0c
44c62006
7c94301c
0016311c
44974664
0007080f
05c31294
1c0ca2d2
c3d216c3
2c0c3ac3
43d228c3
540c5dc3
60376006
0b1ea4bc
04739066
0ebc0457
30c30892
04573364
649713c3
64d74c0c
0ac9dabc
000740c3
05c31454
1c0ca2d2
c3d216c3
340c5ac3
43d228c3
4c0c3dc3
740ca497
a037a006
0b1ea4bc
80060053
019604c3
0f56fc76
00000804
0f36f016
90c3ba96
42c381c3
51774006
0ebc01c3
b0c30892
4006b364
50f75137
40774037
40f740b7
41774137
41f741b7
1f3c04c3
2f3c1140
60061100
0b1f62bc
000750c3
000c74dc
10f8701c
0000711c
8c0c7c0c
0098001c
44c615c3
7c60301c
0016311c
60c34664
14540007
8c0c7c0c
15c31117
301c44c6
311c7c60
46640016
0af270c3
1157a037
25c315c3
a4bc35c3
b0660b1e
af5c13f3
06c30884
f4bc15c3
50c30b1c
600607d2
11576037
23c313c3
931c09b3
20940002
02004f3c
bcbc04c3
04c30b1d
2bc318c3
0b1daabc
0cc09f3c
19c304c3
0b1d9abc
77b8001c
0016011c
10c01f3c
301c26c3
38bc04a8
80c30b1c
16540007
06c30133
0b1ce6bc
1157a037
25c317c3
06c30af3
0b1ce6bc
1157a037
25c317c3
a4bc35c3
58c30b1e
c0370b73
09c3a077
27c32406
86bc3ac3
50c30b1c
23c37117
0d5402e4
e6bc06c3
8f5c0b1c
11570007
28c317c3
a4bc32c3
08530b1e
315707c3
eabc25c3
40c308cb
06c30ad2
0b1ce6bc
00078f5c
17c31157
045328c3
08c08f3c
07c3c037
28c33117
5abc6806
50c30b1c
09540407
e6bc06c3
80370b1c
17c31157
fb3324c3
19c308c3
eabc25c3
0dd208cb
e6bc06c3
40060b1c
11574037
32c317c3
0b1ea4bc
0193bfe6
e6bc06c3
60060b1c
11576037
26c317c3
0b1ea4bc
05c3a006
f0764696
08040f56
b396f016
41c370c3
73376006
08920ebc
636460c3
72f76006
60776037
60f760b7
61776137
61f761b7
1f3c04c3
2f3c1300
62bc12c0
40c30b1f
38940007
02005f3c
8cbc05c3
40c30b1d
05c308f2
26c317c3
0b1d7abc
05d240c3
60376006
01b31317
0ec06f3c
16c305c3
0b1d6abc
331740c3
600607d2
01c36037
23c313c3
06c302b3
eabc4806
331708cb
80370ad2
14c301c3
34c324c3
0b1ea4bc
01139fe6
01c38037
24c314c3
a4bc34c3
04c30b1e
0f564d96
00000804
b796f016
41c370c3
72376006
08920ebc
636460c3
71f76006
60776037
60f760b7
61776137
61f761b7
1f3c04c3
2f3c1200
62bc11c0
40c30b1f
38940007
02005f3c
5cbc05c3
40c30b1d
05c308f2
26c317c3
0b1d4abc
05d240c3
60376006
01b31217
0ec06f3c
16c305c3
0b1d3abc
321740c3
600607d2
01c36037
23c313c3
06c302b3
eabc4606
321708cb
80370ad2
14c301c3
34c324c3
0b1ea4bc
01139fe6
01c38037
24c314c3
a4bc34c3
04c30b1e
0f564996
00000804
d396f016
41c370c3
6b376006
08920ebc
636460c3
6af76006
60776037
60f760b7
61776137
61f761b7
1f3c04c3
2f3c0b00
62bc0ac0
40c30b1f
38940007
02005f3c
bcbc05c3
40c30b1d
05c308f2
26c317c3
0b1daabc
05d240c3
60376006
01b30b17
08c06f3c
16c305c3
0b1d9abc
2b1740c3
600607d2
01c36037
23c313c3
06c302b3
eabc4406
2b1708cb
80370ad2
14c301c3
34c324c3
0b1ea4bc
01139fe6
01c38037
24c314c3
a4bc34c3
04c30b1e
0f562d96
00000804
a496f016
200641c3
36b736f7
36373677
35b735f7
35373577
16801f3c
1f3c2037
20771580
2f3c40b7
40f71640
15402f3c
61774137
16003f3c
3f3c61b7
61f71500
16c01f3c
15c02f3c
62bc34c3
50c30b1f
75940007
10f8301c
0000311c
8c0c6c0c
15c31557
301c44c6
311c7c80
46640016
36d740c3
0af27697
01c3a037
565713c3
a4bc7617
b0660b1e
7f3c0b53
a0370200
55d707c3
0b1e8cbc
565750c3
32940007
14c307c3
68bc7557
50c30b1e
06d2d617
16d78037
56573697
04c307f3
555716c3
08cbeabc
769736d7
803707d2
13c301c3
76175657
40260553
07c34037
8cbc55d7
50c30b1e
803706d2
369716d7
01b35657
14c307c3
755724c3
0b1e54bc
565750c3
803706d2
369716d7
02f37617
12c304c3
eabc5557
36d708cb
56577697
09d2d617
01c38037
36c313c3
0b1ea4bc
00f3bfe6
01c38037
36c313c3
0b1ea4bc
5c9605c3
08040f56
001cfc96
011c6cc0
101c0016
111c6d04
201c0016
211c6d28
301c0016
311c6dcc
94bc0016
00070b22
001c6894
011c6e70
101c0016
111c6e94
201c0016
211c6eb8
301c0016
311c6f3c
94bc0016
00070b22
001c5494
011c6fc0
101c0016
111c6fc4
3abc0016
00070b22
001c4b94
011c6fc0
101c0016
111c7008
e0bc0016
00070b21
001c3f94
011c6fc0
101c0016
111c706c
86bc0016
00070b21
00463394
70f0101c
0016111c
710c201c
0016211c
0b2098bc
28940007
7594301c
0016311c
301c6037
3f5c0200
301c0026
311c7590
60b70016
3f5c6066
001c0066
011c7310
101c0016
201c0080
211c7390
301c0016
d6bc0200
30c30b1e
00d369d2
ff34001c
1fe600b3
001c0073
0496ff31
00000804
1420201c
0000211c
63f2680c
680f6026
08040006
08040006
08040006
08040006
08040006
019e301c
1c5400a7
0bb400a7
13540067
00676b06
301c15b4
0027ff18
02130f94
01a0301c
0c5400e7
019f301c
081400e7
04940107
0289301c
301c0073
03c3ff53
00000804
00a76406
00a71554
620608b4
10540067
00876286
01930b94
00e76806
66060954
061400e7
01076486
301c0354
03c3ff53
00000804
e6bc4b86
080408cb
e6bc4c06
080408cb
e6bc4d86
080408cb
0336f016
81c370c3
301c92c3
311c10f8
6c0c0000
001c8c0c
200600cc
301c44c6
311c7cb0
46640016
b06660c3
1f540007
0b1d5cbc
0df250c3
17c306c3
4abc28c3
50c30b1d
06c306f2
3abc19c3
50c30b1d
10f8301c
0000311c
8c4c6c0c
200606c3
301c44c6
311c7cb0
46640016
c07605c3
08040f56
cd967016
61c350c3
24f202d2
ff53601c
0fc30253
201c15c3
e6bc00cc
05c308cb
3abc16c3
60c30b1d
1fc305c3
00cc201c
08cbe6bc
339606c3
08040e56
0336f016
81c370c3
301c92c3
311c10f8
6c0c0000
001c8c0c
200600cc
301c44c6
311c7cc0
46640016
b06660c3
1f540007
0b1d8cbc
0df250c3
17c306c3
7abc28c3
50c30b1d
06c306f2
6abc19c3
50c30b1d
10f8301c
0000311c
8c4c6c0c
200606c3
301c44c6
311c7cc0
46640016
c07605c3
08040f56
cd967016
61c350c3
24f202d2
ff53601c
0fc30253
201c15c3
e6bc00cc
05c308cb
6abc16c3
60c30b1d
1fc305c3
00cc201c
08cbe6bc
339606c3
08040e56
0336f016
81c370c3
301c92c3
311c10f8
6c0c0000
0d868c0c
44c62006
7cd0301c
0016311c
60c34664
0007b066
bcbc1f54
50c30b1d
06c30df2
28c317c3
0b1daabc
06f250c3
19c306c3
0b1d9abc
301c50c3
311c10f8
6c0c0000
06c38c4c
44c62006
7cd0301c
0016311c
05c34664
0f56c076
00000804
e596f016
51c340c3
0fc3ed86
27c314c3
08cbe6bc
15c304c3
0b1d9abc
04c350c3
27c31fc3
08cbe6bc
1b9605c3
08040f56
0336f016
81c370c3
301c92c3
311c10f8
6c0c0000
0c068c0c
44c62006
7ce0301c
0016311c
50c34664
0007d066
ecbc1c54
60c30b1d
05c30af2
28c317c3
0b1ddabc
19c305c3
0b1dcabc
10f8301c
0000311c
8c4c6c0c
200605c3
301c44c6
311c7ce0
46640016
c07606c3
08040f56
e896f016
51c340c3
0fc3ec06
27c314c3
08cbe6bc
15c304c3
0b1dcabc
04c350c3
27c31fc3
08cbe6bc
189605c3
08040f56
e996f016
71c340c3
0fc3cb86
26c314c3
08cbe6bc
17c304c3
0b055cbc
1fc304c3
e6bc26c3
179608cb
08040f56
40c3f016
62c351c3
f0bc73c3
20c30b23
ff7c001c
32e46157
80a73b14
80a71b54
806706b4
80870d54
02130894
1e5480e7
161480e7
20548107
ff53001c
05c30533
27c316c3
0b05d2bc
05c30473
27c316c3
05c303b3
27c316c3
0b24c6bc
05c30333
27c316c3
0b2416bc
05c30273
27c316c3
0b246ebc
05c301b3
27c316c3
0b05d2bc
05c307f2
273c16c3
18bc0100
0f560b25
00000804
0736f016
80c3ff96
a2c391c3
301c73c3
311c10f8
6c0c0000
001c8c0c
20060130
301c44c6
311c7cec
46640016
b06660c3
1f540007
60376006
425717c3
8cbc6297
50c30b1e
06c308f2
29c318c3
68bc3ac3
50c30b1e
10f8301c
0000311c
8c4c6c0c
200606c3
301c44c6
311c7cec
46640016
019605c3
0f56e076
00000804
0736f016
80c3ff96
a2c391c3
301c73c3
311c10f8
6c0c0000
001c8c0c
20060130
301c44c6
311c7d04
46640016
b06660c3
1f540007
60376026
425717c3
8cbc6297
50c30b1e
06c308f2
29c318c3
54bc3ac3
50c30b1e
10f8301c
0000311c
8c4c6c0c
200606c3
301c44c6
311c7d04
46640016
019605c3
0f56e076
00000804
00000000
00000000
00000000
00000000
415f6377
62437365
636e4563
74707972
00000000
415f6377
6e457365
70797263
00000074
00180005
3d4e432f
00000000
3d4e532f
00000000
003d432f
003d4c2f
3d54532f
00000000
003d4f2f
3d554f2f
00000000
7265732f
4e6c6169
65626d75
00003d72
616d652f
64416c69
73657264
00003d73
4449552f
0000003d
2d2d2d2d
4745422d
43204e49
49545245
41434946
2d2d4554
002d2d2d
2d2d2d2d
444e452d
52454320
49464954
45544143
2d2d2d2d
0000002d
2d2d2d2d
4745422d
43204e49
49545245
41434946
52204554
45555145
2d2d5453
002d2d2d
2d2d2d2d
444e452d
52454320
49464954
45544143
51455220
54534555
2d2d2d2d
0000002d
2d2d2d2d
4745422d
44204e49
41502048
454d4152
53524554
2d2d2d2d
0000002d
2d2d2d2d
444e452d
20484420
41524150
4554454d
2d2d5352
002d2d2d
2d2d2d2d
4745422d
58204e49
20393035
2d4c5243
2d2d2d2d
00000000
2d2d2d2d
444e452d
30355820
52432039
2d2d2d4c
00002d2d
2d2d2d2d
4745422d
52204e49
50204153
41564952
4b204554
2d2d5945
002d2d2d
2d2d2d2d
444e452d
41535220
49525020
45544156
59454b20
2d2d2d2d
0000002d
2d2d2d2d
4745422d
50204e49
41564952
4b204554
2d2d5945
002d2d2d
2d2d2d2d
444e452d
49525020
45544156
59454b20
2d2d2d2d
0000002d
2d2d2d2d
4745422d
45204e49
5952434e
44455450
49525020
45544156
59454b20
2d2d2d2d
0000002d
2d2d2d2d
444e452d
434e4520
54505952
50204445
41564952
4b204554
2d2d5945
002d2d2d
2d2d2d2d
4745422d
45204e49
52502043
54415649
454b2045
2d2d2d59
00002d2d
2d2d2d2d
444e452d
20434520
56495250
20455441
2d59454b
2d2d2d2d
00000000
2d2d2d2d
4745422d
44204e49
50204153
41564952
4b204554
2d2d5945
002d2d2d
2d2d2d2d
444e452d
41534420
49525020
45544156
59454b20
2d2d2d2d
0000002d
2d2d2d2d
4745422d
50204e49
494c4255
454b2043
2d2d2d59
00002d2d
2d2d2d2d
444e452d
42555020
2043494c
2d59454b
2d2d2d2d
00000000
65657246
7073634f
75716552
00747365
74696e49
7073634f
75716552
00747365
0501062b
01300705
00000002
666e6f43
536d7269
616e6769
65727574
00000000
455f6377
72506363
74617669
79654b65
6f636544
00006564
65657246
6e676953
00007265
656b614d
6e676953
00007265
6f636544
6c416564
6d614e74
00007365
6f636544
75536564
65727462
00000065
73726150
72654365
00000074
8648862a
02020df7
8648862a
05020df7
02030e2b
0000001a
01488660
02040365
00000001
01488660
02040365
00000002
01488660
02040365
00000003
ce48862a
00030438
8648862a
01010df7
00000002
8648862a
01010df7
00000004
8648862a
01010df7
00000005
8648862a
01010df7
0000000b
8648862a
01010df7
0000000c
8648862a
01010df7
0000000d
ce48862a
0001043d
ce48862a
0203043d
ce48862a
0303043d
ce48862a
0403043d
ce48862a
00010438
8648862a
01010df7
00000001
ce48862a
0001023d
02030e2b
00000007
8648862a
07030df7
0501062b
01300705
00000001
0501062b
01300705
00000002
00131d55
00111d55
001f1d55
0501062b
01010705
00231d55
000e1d55
00201d55
000f1d55
00361d55
00251d55
001e1d55
0501062b
01300705
0501062b
02300705
00201d55
0501062b
04080705
00251d55
0501062b
01030705
0501062b
02030705
0501062b
09030705
8648862a
05010df7
0000000c
4e746547
00656d61
4b746547
00007965
65657246
6f636544
43646564
00747265
65657246
656d614e
74627553
73656572
00000000
65657246
4e746c41
73656d61
00000000
72546f54
74696461
616e6f69
636e456c
00000000
72636544
4b747079
00007965
03020100
07060504
ffff0908
ffffffff
0c0b0aff
ff0f0e0d
ffffffff
ffffffff
ffffffff
ffffffff
ffffffff
ffffffff
0c0b0aff
000f0e0d
44434241
48474645
4c4b4a49
504f4e4d
54535251
58575655
62615a59
66656463
6a696867
6e6d6c6b
7271706f
76757473
7a797877
33323130
37363534
2f2b3938
ffffff3e
3635343f
3a393837
ff3d3c3b
ffffffff
0100ffff
05040302
09080706
0d0c0b0a
11100f0e
15141312
19181716
ffffffff
1b1affff
1f1e1d1c
23222120
27262524
2b2a2928
2f2e2d2c
33323130
50434553
52323131
00000031
43374244
46424132
33453236
36364535
36373038
44414542
42383032
00000000
43374244
46424132
33453236
36364535
36373038
44414542
38383032
00000000
45393536
41423846
39333430
45453631
39384544
30373131
32324232
00000000
43374244
46424132
33453236
36374535
46443832
35364341
35433136
00000000
37383439
39393332
35413539
36374545
46353542
46324339
00383930
43393841
46413545
34323738
32413043
45304533
37464630
30303537
00000000
50434553
52383231
00000031
46464646
44464646
46464646
46464646
46464646
46464646
46464646
46464646
00000000
46464646
44464646
46464646
46464646
46464646
46464646
46464646
43464646
00000000
35373845
31433937
39373031
44333446
34323844
43333939
45454332
33444535
00000000
46464646
45464646
30303030
30303030
33413537
42314430
38333039
35313141
00000000
46313631
32353746
39384238
44324239
38324330
43373036
43323541
36384235
00000000
41354643
39333843
46414235
33314245
44323043
32393241
44454444
33384137
00000000
50434553
52303631
00000031
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464637
46464646
00000000
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464637
43464646
00000000
37394331
43464542
44423435
42384137
43413536
46393846
34443138
44413444
35363543
35344146
00000000
30303031
30303030
30303030
30303030
30303030
43344631
32394638
44454137
37414333
35323235
00000037
36394134
38363542
35464538
38323337
34363634
39383936
33433836
39424238
42433331
32384346
00000000
36413332
35353832
38363133
44373439
43443935
32313943
33323430
37333135
35434137
32334246
00000000
50434553
52323931
00000031
46464646
46464646
46464646
46464646
46464646
46464646
46464646
45464646
46464646
46464646
46464646
46464646
00000000
46464646
46464646
46464646
46464646
46464646
46464646
46464646
45464646
46464646
46464646
46464646
43464646
00000000
31323436
39313530
43393545
37453038
37414630
42413945
34323237
39343033
38424546
43454544
36343143
31423942
00000000
46464646
46464646
46464646
46464646
46464646
46464646
45443939
36333846
42363431
31423943
32443442
31333832
00000000
44383831
45303841
30333042
36463039
46424337
42453032
31413334
30303838
46463446
44464130
46463238
32313031
00000000
32393137
46353942
44384346
36383741
31303133
36444531
43343242
37354444
37394633
31314137
34393745
00313138
50434553
52343232
00000031
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
30303030
30303030
30303030
30303030
30303030
31303030
00000000
46464646
46464646
46464646
46464646
46464646
46464646
46464646
45464646
46464646
46464646
46464646
46464646
46464646
45464646
00000000
35303442
35384130
34304330
42413342
31343546
36353233
34343035
37423042
46423744
41423844
42303732
33343933
35353332
34424646
00000000
46464646
46464646
46464646
46464646
46464646
46464646
46464646
32413631
38423045
45333046
44443331
35343932
43354335
44334132
00000000
45303742
44424330
34424236
46374642
33313233
39423039
33304134
33443143
32433635
32323131
32333433
36443038
43353131
31324431
00000000
37334442
38383336
37463542
42463332
32324334
36454644
33344443
30413537
37304135
34363734
35443434
39393138
30303538
34334537
00000000
4d495250
39333245
00003156
46464637
46464646
46464646
46464646
46464646
46464646
46464637
46464646
46464646
30303038
30303030
30303030
46464637
46464646
46464646
00000000
46464637
46464646
46464646
46464646
46464646
46464646
46464637
46464646
46464646
30303038
30303030
30303030
46464637
46464646
43464646
00000000
31304236
42334336
31464344
31343938
36443044
32393435
35373431
31374143
42443941
32424632
44314437
39373733
35383136
34393243
41304332
00000000
46464637
46464646
46464646
46464646
46464646
46464646
46464637
45394646
41394535
44354639
31373039
31444246
36323235
30393838
42304439
00000000
41464630
43333639
38414344
43363138
33334343
34363842
44454232
35303946
33443343
37353835
46334433
42463732
42334442
39424333
46414141
00000000
42454437
34453845
41303945
45414435
30344536
41433435
42303335
36343041
33423435
38313836
32324543
39334236
42434346
32304237
45413146
00000000
50434553
52363532
00000031
46464646
46464646
30303030
31303030
30303030
30303030
30303030
30303030
30303030
30303030
46464646
46464646
46464646
46464646
46464646
46464646
00000000
46464646
46464646
30303030
31303030
30303030
30303030
30303030
30303030
30303030
30303030
46464646
46464646
46464646
46464646
46464646
43464646
00000000
36434135
38443533
41334141
37453339
42453342
35354442
38393637
43423638
44313536
30423630
33354343
36463042
45434233
45334333
32443732
42343036
00000000
46464646
46464646
30303030
30303030
46464646
46464646
46464646
46464646
36454342
44414146
37313741
34384539
39423346
32434143
33364346
31353532
00000000
37314236
32463144
43323145
37343234
43423846
35453645
34413336
32463034
33303737
31384437
42454432
30413333
31413446
35343933
38393844
36393243
00000000
33454634
32453234
41314546
42394637
37454538
41344245
46304337
36314539
45434232
37353333
31334236
45434535
36424243
38363034
46423733
35463135
00000000
50434553
52343833
00000031
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
45464646
46464646
46464646
30303030
30303030
30303030
30303030
46464646
46464646
00000000
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
45464646
46464646
46464646
30303030
30303030
30303030
30303030
46464646
43464646
00000000
31333342
37414632
45333245
34453745
45383839
42363530
38463345
39314432
44313831
45364339
31384546
32313134
34313330
46383830
33313035
41353738
36353643
44383933
45324138
44393144
35384132
44453843
43453344
46454132
00000000
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
33363743
31384434
37333446
46444432
41313835
32424430
30423834
41373741
43454345
41363931
35434343
33373932
00000000
37384141
32324143
42384542
37333530
31424538
45313743
30323346
34374441
44314536
32364233
37414238
38394239
37463935
30453134
34353238
38334132
32303535
44353246
35354642
43363932
34354133
38334535
36373237
37424130
00000000
37313633
41344544
36323639
46364332
45394435
46423839
32393239
39324344
34463846
44424431
41393832
43373431
41443945
33313133
30463542
30433842
30364130
45433142
45374431
44393138
33344137
43374431
41453039
46354530
00000000
50434553
52313235
00000031
46464631
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
00464646
46464631
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
00434646
35393135
39424533
45383136
41394331
32394631
31324139
36423041
30343538
32414545
32374144
39394235
35313342
38423346
39383442
45383139
39303146
36353145
39333931
43453135
33394537
36314237
30433235
42334442
46423142
35333730
46443337
44333838
34334332
46453146
46313534
42363444
46333035
00003030
46464631
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
46464646
35414646
38363831
42333837
39463246
37423636
30434346
46383431
41393037
33304435
43354242
38384239
34433939
42454137
42463642
39453137
36383331
00393034
35383643
36304538
34303742
39453430
45394443
42434533
33323636
34423539
43393234
31383436
35303933
35424633
38463132
46413832
42363036
44334434
31414142
45354234
46453737
39353745
45463832
31434431
32413732
38414646
33334544
33423834
35383143
32344136
39464239
45374537
32433133
44423545
00003636
33383131
36393239
39383741
43423341
35343030
35413843
32344246
31443743
39394442
34354638
35393434
34423937
31383634
42464137
32373144
36453337
39433236
37454537
35393932
32344645
43303436
42303535
33313039
30444146
33313637
37433335
41363830
43323732
38303432
39454238
39363734
36314446
00303536
0000000e
00000008
001652a8
001652b4
001652d4
001652f4
00165314
00165334
00165350
00166344
00000005
000000b6
00000001
00000010
0000000a
00165370
0016537c
001653a0
001653c4
001653e8
0016540c
00165430
0016634c
00000005
000000cc
00000001
00000014
0000000c
00165454
00165460
0016548c
001654b8
001654e4
00165510
0016553c
00166354
00000005
000000b8
00000001
00000018
00000001
00165568
00165574
001655a8
001655dc
00165610
00165644
00165678
0016635c
00000008
00000208
00000001
0000001c
0000000e
001656a8
001656b4
001656f0
0016572c
00165768
001657a4
001657e0
00166364
00000005
000000d1
00000001
0000001e
00000004
0016581c
00165828
00165868
001658a8
001658e8
00165928
00165968
0016636c
00000008
0000020b
00000001
00000020
00000007
001659a8
001659b4
001659f8
00165a3c
00165a80
00165ac4
00165b08
00166374
00000008
0000020e
00000001
00000030
0000000f
00165b4c
00165b58
00165bbc
00165c20
00165c84
00165ce8
00165d4c
0016637c
00000005
000000d2
00000001
00000042
00000010
00165db0
00165dbc
00165e40
00165ec4
00165f48
00165fcc
00166050
00166384
00000005
000000d3
00000001
00000000
ffffffff
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
655f6377
655f6363
726f7078
39785f74
00003336
655f6377
655f6363
726f7078
6f705f74
5f746e69
00726564
655f6377
6d5f6363
5f656b61
5f79656b
00007865
655f6377
645f6363
705f6c65
746e696f
0000685f
655f6377
6e5f6363
705f7765
746e696f
0000685f
0004812b
00000006
0004812b
0000001c
0004812b
00000008
ce48862a
0101033d
0004812b
00000021
ce48862a
0401033d
ce48862a
0701033d
0004812b
00000022
0004812b
00000023
485f6377
0046444b
00180005
001667a0
001667a0
00000002
00000003
00000005
00000007
0000000b
0000000d
00000011
00000013
00000017
0000001d
0000001f
00000025
00000029
0000002b
0000002f
00000035
0000003b
0000003d
00000043
00000047
00000049
0000004f
00000053
00000059
00000061
00000065
00000067
0000006b
0000006d
00000071
0000007f
00000083
00000089
0000008b
00000095
00000097
0000009d
000000a3
000000a7
000000ad
000000b3
000000b5
000000bf
000000c1
000000c5
000000c7
000000d3
000000df
000000e3
000000e5
000000e9
000000ef
000000f1
000000fb
00000101
00000107
0000010d
0000010f
00000115
00000119
0000011b
00000125
00000133
00000137
00000139
0000013d
0000014b
00000151
0000015b
0000015d
00000161
00000167
0000016f
00000175
0000017b
0000017f
00000185
0000018d
00000191
00000199
000001a3
000001a5
000001af
000001b1
000001b7
000001bb
000001c1
000001c9
000001cd
000001cf
000001d3
000001df
000001e7
000001eb
000001f3
000001f7
000001fd
00000209
0000020b
0000021d
00000223
0000022d
00000233
00000239
0000023b
00000241
0000024b
00000251
00000257
00000259
0000025f
00000265
00000269
0000026b
00000277
00000281
00000283
00000287
0000028d
00000293
00000295
000002a1
000002a5
000002ab
000002b3
000002bd
000002c5
000002cf
000002d7
000002dd
000002e3
000002e7
000002ef
000002f5
000002f9
00000301
00000305
00000313
0000031d
00000329
0000032b
00000335
00000337
0000033b
0000033d
00000347
00000355
00000359
0000035b
0000035f
0000036d
00000371
00000373
00000377
0000038b
0000038f
00000397
000003a1
000003a9
000003ad
000003b3
000003b9
000003c7
000003cb
000003d1
000003d7
000003df
000003e5
000003f1
000003f5
000003fb
000003fd
00000407
00000409
0000040f
00000419
0000041b
00000425
00000427
0000042d
0000043f
00000443
00000445
00000449
0000044f
00000455
0000045d
00000463
00000469
0000047f
00000481
0000048b
00000493
0000049d
000004a3
000004a9
000004b1
000004bd
000004c1
000004c7
000004cd
000004cf
000004d5
000004e1
000004eb
000004fd
000004ff
00000503
00000509
0000050b
00000511
00000515
00000517
0000051b
00000527
00000529
0000052f
00000551
00000557
0000055d
00000565
00000577
00000581
0000058f
00000593
00000595
00000599
0000059f
000005a7
000005ab
000005ad
000005b3
000005bf
000005c9
000005cb
000005cf
000005d1
000005d5
000005db
000005e7
000005f3
000005fb
00000607
0000060d
00000611
00000617
0000061f
00000623
0000062b
0000062f
0000063d
00000641
00000647
00000649
0000064d
00000653
00000004
00000000
00000001
00000000
00000002
00000000
00000001
00000000
00000003
00000000
00000001
00000000
00000002
00000000
00000001
00000000
74736166
6d5f735f
756d5f70
69685f6c
645f6867
00736769
74736166
6d5f735f
756d5f70
69645f6c
00007367
74736166
6d5f735f
71735f70
00000072
695f706d
5f74696e
657a6973
00000000
74736166
5f706d5f
746e6f6d
656d6f67
725f7972
63756465
00000065
675f706d
00776f72
665f706d
6563726f
6f72657a
00000000
635f706d
7261656c
00000000
695f706d
0074696e
33323130
37363534
42413938
46454443
4a494847
4e4d4c4b
5251504f
56555453
5a595857
64636261
68676665
6c6b6a69
706f6e6d
74737271
78777675
2f2b7a79
00000000
4835644d
00687361
505f6377
3153434b
42505f32
5f46444b
00007865
505f6377
46444b42
00000032
f3d05aa6
0e4edb45
c375e8ff
421fe7a2
629d12c7
19c1f50f
f055efa9
fbe08551
31f98185
6e271775
7d60e906
2ecccbdb
77333663
46861ee4
b40aeb8d
3f68eda8
474e136a
00c714e0
e9814e45
69a55853
8fa38a80
23a6722a
9f5a9159
68ca048a
8e8a2be6
b641f1e8
e3660598
49c0e3bf
acd4da03
229fdf2c
670a0180
d383bc39
e38f2f6e
4289cdcd
0b8919bc
d39de870
fb6df47e
09c217dc
231b1b94
70b31764
bbe5e24a
009528bf
5bd48f06
9cb6406b
614f9478
00cf5512
50ee5f66
04c6d7d6
19686df9
50afbf2e
198aa88e
cd9c7b3c
3470a404
a9e57dee
9b709a54
8bb30172
e8df7f30
e81bff42
e6bcfcf7
00282ac8
5d60ab32
51568ddc
598a3b09
de3a9dbd
219e24a1
4a2e9ea6
5f516739
1cd43aa0
6e125bcf
68b2f3b9
2d950c08
fe4182f8
bc7bc24c
00d5bebb
1d69a28e
b4eb1519
ca935597
bad0ba3f
d9267013
5059a901
1dc407a2
153e77c7
4a5fe8c1
2800915f
eb0b8366
17eec4e5
3239b885
0044bb3f
937d1759
50053f84
a53339f3
1688b41e
9cab9986
36156585
c77e1fa6
4a278b1e
e5171f15
53afec6b
55c9cf1d
b6adf1f2
b2516d53
003cd556
69027c89
e154429f
f7943cf3
a35da8bf
c2f66d82
81d00e59
36edbc5c
37a37ad7
ff82155a
4187c8c1
a01bfd6a
df6d4bf0
0e2b1af8
004d845b
77333663
46861ee4
b40aeb8d
3f68eda8
474e136a
00c714e0
e9814e45
69a55853
8fa38a80
23a6722a
9f5a9159
68ca048a
8e8a2be6
b641f1e8
e3660598
49c0e3bf
acd4da03
229fdf2c
670a0180
d383bc39
3bc6ee04
2cdf31b2
fb1a0a63
9d9424e7
78585a00
79aae151
4773475e
6256b0c8
dcbd181c
fc998ddd
20b9c25f
accfd853
83b80bfb
d1fa0512
71c0d6dd
18608a31
f5733bf0
d0d4e4ed
03def971
10ea7afd
b899925d
07aa99af
b94ddb5b
8dc128aa
ee564b17
094d012a
22ff9688
a855c982
69e06919
07e08cfa
3a1880a1
17aedf07
f3d05aa6
0e4edb45
c375e8ff
421fe7a2
629d12c7
19c1f50f
f055efa9
fbe08551
31f98185
6e271775
7d60e906
2ecccbdb
c360e1d3
40f3995b
648262b2
601075d1
a35d04e0
a557ff83
73a6737d
0dd8b8d2
c3a6f6aa
45bb915a
d03fd779
11d1fec8
061339b0
eddf8a82
81018f52
bdfeb321
97e743c3
63bb7db8
de3313db
e1ecd1d9
b7a6cf77
1dabe81f
ed2466a4
1ce51564
cac7e2cd
9983e286
91ebea0e
52150412
9195228b
2db08102
c9f431d4
df2704f7
525f6377
485f474e
746c6165
73655468
00000074
465f6377
52656572
0000676e
525f6377
485f474e
746c6165
73655468
636f4c74
00006c61
495f6377
5274696e
655f676e
00000078
50617352
4f5f6461
00504541
4d617352
00314647
50617352
61766972
65446574
70797263
00784574
55617352
6461506e
45414f5f
00000050
525f6377
6c436173
756e6165
00000070
62386539
66633637
30646265
32323136
32303166
62343434
31306533
66333364
64383363
38656131
66663339
37373236
36333865
63663835
35643736
33336336
00000000
35623233
34343836
66333463
34356334
63636539
63306638
37313333
35313464
00000000
66313831
62653736
63656166
34663765
39613238
64333566
31303039
31376339
33613262
38343665
30613035
39306161
34313632
64343661
39303766
35306463
38393038
65623265
31356361
34323634
65643630
35636630
32653337
38313935
37323132
65623165
39666262
37303064
64636664
38623464
37323164
63303537
61623137
38663761
30646136
33626239
63656461
36376264
65616531
31383639
00000000
66663532
64313438
38613865
63306234
65653966
61303239
34366231
34653934
37616439
34366663
34633262
34656234
34373230
32363466
32663964
61653734
39656239
63303031
66326331
64623466
62626231
39636136
30636238
64386632
64336166
31393765
39663661
34373364
65646136
39373963
66316165
31323566
35346634
61333738
62363839
38633633
61383533
39646137
36663365
33326464
00000000
65376232
36313531
65613832
36613264
37666261
38383531
66633930
63336634
00000000
31303030
33303230
35303430
37303630
39303830
62306130
64306330
66306530
00000000
31636236
32656562
30346532
36396639
64333965
31316537
33393337
61323731
64326561
37356138
33306531
63396361
37626539
63616636
66613534
31356538
38633033
36346331
63353361
31313465
62663565
39313163
61306131
66653235
66393666
35343432
66346664
37316239
62326461
62373134
63363665
30313733
00000000
39343637
63616261
39313138
36343262
39656563
62396538
39653231
64373931
36383035
62396263
32373035
65653931
62643539
61333131
36373139
32623837
65623337
38623664
31633365
62333437
36313137
65393665
32323232
36313539
31666633
31616163
66313836
39306361
65303231
30336163
36383537
37613165
00000000
00636261
38376162
66623631
31306638
61656663
31343134
65643034
65616435
33323232
33303062
33613136
37313639
63396137
30313462
31366666
30303266
64613531
00000000
30306263
66333537
33613534
62386535
30613562
39366433
36636139
37303035
63323732
62613233
65646530
33363164
62386131
61353036
66663334
64656235
36383038
62323730
37653161
33326363
61623835
31616365
38633433
37613532
00000000
66616464
31613533
31363339
61626137
31346363
39343337
30326561
31333134
36653231
65346166
39613938
32616537
65396130
36656565
35356234
61393364
32393132
61323939
66343732
38613163
61623633
33326333
65663361
64626265
64343534
33323434
63333436
65303865
61396132
66343963
63343561
66393461
00000000
72657645
656e6f79
74656720
72462073
79616469
66666f20
0000002e
41464338
37393735
38373539
37443942
37433138
45453746
31324444
32363945
35344346
37423844
41444343
33383836
34384437
34333845
33373935
30363538
30433938
30413532
39384636
44373746
36334337
34433439
36413338
42364645
45453234
38423936
30453243
31434331
31463331
34463733
39383839
32353730
43364645
34393036
31383344
39373939
37323231
45383239
44323844
35424235
39424630
35374136
37394634
36364437
35374546
46434241
35463037
34343944
32353338
33443632
36464230
44323646
43394237
41464641
37313831
44354339
45434241
41423835
34373934
35413432
44384341
38313136
37423431
46433632
34393233
32433044
30303833
32434430
35373742
39313937
41433532
46383235
39344236
33443734
41423445
43384631
43344644
38384533
41413145
44434632
36344541
44364631
35343246
43334444
39463933
44463038
43454630
46333132
42374243
36314437
34463937
44393836
33353830
36314538
30453841
37353346
46444142
30463144
43363544
42353336
45364539
44424337
46324536
33463233
42413734
37304539
31353836
31303636
46454536
35384638
35373337
38313234
35333635
34383836
43423936
46413830
42333437
35423230
42463643
44454335
34323938
43303242
42373431
34334639
41414639
33343931
36464244
41433737
00000000
61eac542
19f0257a
72e19e32
852493e4
d0ab8d51
91248319
73745989
6c61a6b4
e68ebac5
1dade093
c8f0e076
fbc0c85a
4cb2ec11
35b72cee
b993758f
4a908bfa
eb7305ec
92af996d
d0d999a8
b35cbefa
ec6e2549
2d429797
d57f0dd6
cff273fe
b77fad5e
3f5ed82f
d284d26f
775efced
f7c53ea0
422f4c3c
0f222807
c3efe9e9
f1df3668
9141a5be
e2cc9c6b
1f925e69
7a737af2
5c4a4fc5
eeac2f3b
3bdda880
936ce8bf
a58dafa1
2ca9b3c6
c7fa5d44
9ffa15e2
58c9673d
8a85ba9d
6a323f22
d0f5b8fe
ac282ff9
c271364e
0b4e5b2b
76f76642
bb28a9ac
9f920903
622b452c
5c6762d4
8e3809ef
0ccf2057
d45193b9
07795940
ce82db20
797e4d01
32832658
0542bd84
30134ec6
ff090ee3
2cf62062
7a113c01
86424fce
26e546cd
5a92c494
27a512ba
91de478e
20d8cd0d
e5eb6f39
6cbc9b17
18accdce
8540bd83
2ee9bd30
b29dc493
2eb4fbc6
97f20597
213b7603
892417a8
891883d2
050506bb
e6400904
b95c7c0f
c32783f5
7ecff7d3
e860ad18
52b6ed77
d499a622
58b3dcac
1e7ec8fb
cf681446
cda882dc
2ef8b17f
37873705
1a74aaf4
03f6dd63
aae1239b
704ed919
99589187
8add5a68
4af6a88d
e07b7093
8e4c35b6
c7ef8a9a
5cb44b48
49cabed0
ef0a4a3a
e8aa6a0b
906b8601
82c58356
ccf939bf
80d86807
31b3e4c6
6b5086da
0c188c29
5ea45ff9
c5832453
14374455
4e8b0868
97378f37
097e396c
f08190f8
baf4b6f0
9992e63b
145ff557
eb6b8fa8
e6706b45
7e22c6fb
a4e8c198
c934f7a6
ed130c08
34fbbc58
21bccb56
50835376
5649f500
07d439d8
a4d87135
4d29a22f
e847a7f1
163af58a
203418df
cdcc0930
4730616d
b92a8739
449ae72b
bc5e1262
9c90ba8b
1bd9b4a2
6c0d529e
922f1c68
6e150f07
5187a631
1d3e9922
6835fc94
00010001
653509b1
a2c15407
eef9547e
04775c52
6b051a5d
1b8cdcae
663d5aa0
2e8e2c32
a09c6841
c56e8e2b
cd31335d
1b164e71
3174c735
41c64015
30b1c30c
32ec5ce6
f1cc7753
05775d8a
37a7fa4a
66685be6
7f622723
df92105d
608bc098
5967baa3
9806149b
2815446f
d6f5f1d2
b8c65efe
bd7d79aa
762816b3
239882b0
701cf87a
76358604
dd2d57af
cf87c466
0f2da832
f860e29f
131668f2
55ec8a20
f5223672
bdb33c0d
6d22b133
a29e5b5b
592c7ac9
53314e05
2fec4968
c097250f
dd21e677
dd220aea
25f91dfb
1c94f1c9
ceaf31d4
8ed29803
abfe6c73
62f0d73d
4c2a5aa6
f3a1dc1d
b403fa2a
7c8bfddd
cec00ca4
2922d42e
3cf053d7
dcbcd8c6
c2b76aa7
da5d3c70
bfa98ad0
0a74279a
8c16238b
7b91556b
c0c1d5d3
1e4dc357
da1114fb
5574ab51
b992bd19
8fea2f43
709acbad
dc3adce5
331d08d3
7b7b5033
e9868899
28662988
e66572dd
7755ab4e
c46c5512
157f3792
b6dc78a0
f0e7a620
87fba151
a3dcef54
d03d25de
5b20d4aa
e4592603
7f30fba4
e3bd4f07
592b7040
47b3ac11
4683d737
c72acf00
3cf8627f
8fa79bcc
1b0211f9
bfd18a9f
ae301442
6991640d
5404b544
63620f2c
235e8ec4
9d86f13e
ccc2eff1
5ea9f4f6
7bdeb24d
92a9b14c
3557f6be
bfb4ba11
728ed52c
f535c2a0
2d18fc6d
b6ffdff4
67a53394
5df31574
5f12f584
57eb0052
6bce8c86
3483c574
310e9917
23c97283
a1dc369a
0988b2a0
34617352
53363930
566e6769
31767265
6e4b5f35
416e776f
6577736e
73655472
00000074
a4048230
02000102
00010182
2bd103c3
32a439fe
c8533b45
7c2a2b84
aabd9a74
4707522a
b236a6d6
d08e3207
c67b69ba
d49e44c3
2dfd4881
678ba268
c875a1bb
d24a2c36
ba8bf71b
eff90dcf
1e81f1ec
47039b7b
cc65bf9a
6924657f
8914e8a6
f734e45b
9314b0c5
3a7b67f5
01e1787a
a6915656
d28d4213
4c9c403c
df86d1ef
0c1b5137
f1f53ba1
e4354aa3
df96cee1
4ebf7e1b
e810d097
813008a8
430b20af
6774c514
6f8232b4
88c2868d
83369940
72401eba
52d71722
b0732465
cd19efce
6c78ffae
0312c07b
0d724ed4
a33b6d50
5e99a33b
0cd9c89d
8ad9b385
db2654d9
bbacfa6d
c44c25ff
71f479d1
184086d3
b563b013
c4304e72
2d868497
15d72f56
aec07ff7
e55bfcf5
d3baa1fb
00010302
01820201
e6a20001
71105fd8
2e9e0864
1e6dd16d
b10ad285
2cce478c
12a06a51
91de539e
ea6d1d4c
77f27b59
d9c6d9aa
e1d8ab8a
2663e416
136cb5ff
a5e3b859
2e1772c8
e56f9f0c
6f763f59
c211b149
29162e5a
8eb7de0d
a2d540dc
a11ee0ee
db97bef4
14966386
600998cd
9c76302d
88e6cd3c
799247ee
e2005a0b
7c115f5e
b708f97d
2a890620
ab00fd5d
b3f0e122
5ea924bc
001f0e26
9a21fe2d
d36d5b53
8294ab2b
d8364368
22c62ff6
5d41b5fc
ea60330d
e87e7da4
5691554b
8f575cd3
2f17941f
9ee9deaa
8acff4a8
e4a08e4c
cfb27356
69c5864f
2024f33c
0c965c8b
3b126bfa
dfc1679a
a5b296c6
9b0d92d5
24684209
50d44510
483917e4
948b35d0
8fde116d
810259ca
24ea0081
3369f9a7
52dc71e9
2821887d
bade492f
cce91672
0d887a47
58845794
b0813a16
a6cfa23f
06b01e6c
e78f0029
dbac7677
5ed9c7ca
90263f9b
38fcae52
bb140090
94580fb4
7e6a2fe7
21414f1c
1f5931d4
8d1a8a4e
226c57a7
7ef4e5d8
cb10a632
0355a564
0527a687
b6d7c38c
ba4db227
8f47da30
8b3dd354
98948d84
8102a558
38d50081
c58fc31b
0b470c93
c592356f
c8468db0
f58f1892
eff70a80
b980fea1
caba2ab5
a55db018
8d93d007
1c049cd8
a68e62d4
ff018126
632a8ace
aa403534
89de806d
4d576a23
93ad6e9e
0b90564e
8b739d6d
3d27ae0c
aaf04ede
67786cc5
9c52946c
2d6c6737
dfafbbef
c43c90a6
968dcf47
b4a9989e
50a6c59f
fbf0b3dc
81021774
09835e80
7cbabd62
7442bfa2
d21c7cf5
0d04c969
3d3e7e85
18c31224
f329f37b
6c760e5f
41e47559
329d6984
ab22cdf3
4aba35b0
d9e53cb2
4f62b658
9ee5de5d
b253ca0a
b39ef72c
795b0a6b
916eec65
f620924e
ed16fcfc
e20c76d3
69b27fec
0e786b13
b464465a
a025b75e
4b3a755a
3e3cc7ef
b826fdf7
0a99c420
c3be739a
81810219
9344ba00
1934ac14
60915f3b
d6b4f7ac
51360581
65e83d53
dc2eafdc
7dc93e61
f0877fb8
82039b3b
72ce3729
b1d5114e
a0070cc1
8d4a9199
cf79ec7f
e9b539f1
f762ec85
64bc7dda
0e3c224d
f551d6f2
c099d887
0f5d2011
e25bfd29
d91cd9ae
fc6d5621
ed5fd084
181c1510
3dc4e721
9ed0d74b
22cf956a
9e7b03c9
fc0160e3
8081022f
cf4bd011
9fb9671b
86477510
c231ae65
59ac30c6
0fd95006
f70670b5
62c8d3f0
6edaa87c
d33f21f6
8aea5f7f
2ad93fab
d251f35e
e33730c2
0d75a32d
34214d1e
5c7057d5
ec72bf89
d5686e4a
337418cd
453a8c4e
4096e68f
19f963eb
dd513a86
f3b04b89
285d9ff9
35be3895
e75ccaab
a1345393
39135d45
a1464265
bff5cd9f
53617352
506e6769
3153434b
5f353176
776f6e4b
736e416e
54726577
00747365
4b736541
6e776f6e
77736e41
65547265
00007473
766e6f43
48747265
6f547865
006e6942
65657246
736e6942
00000000
535f6377
38336168
73614834
00000068
535f6377
31356168
73614832
00000068
535f6377
35326168
73614836
00000068
535f6377
61486168
00006873
415f6377
62437365
636e4563
74707972
68746957
0079654b
415f6377
62437365
63654463
74707972
68746957
0079654b
0014a624
0014a61c
0014a614
0014eb34
0016466c
00174e1c
0014a1a4
0014a008
0014a3fc
00149ef4
00149e20
0010fb0c
0010f8a8
0010f978
0010f910
0010f958
0010f288
0010f534
0010f788
0010f190
0014e748
0014e748
0014ed0c
0014e6ec
01c330c3
023513e4
080403c3
305c10c3
00061561
08946067
1569215c
0b0d323c
7f3233c4
080403c3
205c30c3
40671561
00060794
1569335c
0d356047
00060173
00fe231c
00060894
1569335c
00fd331c
002602b4
00000804
1e01005c
00000804
1e24305c
0b8b033c
00000804
00b7fd96
503220c3
2f5c4077
440d0021
48324097
2f5c4037
442d0001
00412f5c
0396444d
00000804
0364fe96
20c30077
40374832
00012f5c
2f5c440d
442d0021
08040296
00f7fc96
583220c3
2f5c40b7
440d0041
503240d7
2f5c4077
442d0021
483240d7
2f5c4037
444d0001
00612f5c
0496446d
00000804
30c31016
40c30049
203c0c09
8c29822c
412c343c
0856640f
00000804
40291016
400942c3
422c323c
0856640e
00000804
30c31016
40c30069
203c0c09
8c29c22c
812c243c
303c0c49
640f412c
08040856
21c3ff96
20372409
202d2829
00012f5c
2026400d
4006204d
0196406d
00000804
422f4006
424f42af
426f42cf
205c42ef
205c0285
08040305
40c3f016
10f8601c
0000611c
701c780c
711c6700
ac4c0017
312c022c
37c343e6
780c5664
12acac4c
43e6312c
566437c3
ac4c780c
312c124c
37c343e6
780c5664
12ccac4c
43e6312c
566437c3
ac4c780c
312c126c
37c343e6
780c5664
12ecac4c
43e6312c
566437c3
08040f56
610d7fe6
614d612d
618d616d
61ad6006
600661ed
602e600e
0804604e
42c33016
21c353c3
18542007
105c20c6
60660985
098d305c
105c20a6
305c0995
6086099d
09a5305c
105c2066
604609ad
09b5305c
09bd105c
80074106
61002954
135c20c6
40250985
20266100
0985135c
61004025
135c20a6
40250985
20266100
0985135c
61004025
135c2086
40250985
20266100
0985135c
61004025
135c2046
40250985
20266100
0985135c
abd24025
20466100
0985135c
61004025
135c2006
40250985
0c56402e
00000804
3f36f016
31c3fc96
436442c3
01e39f5c
02231f5c
6f5c20b7
1f5c0243
4c290263
b01c6c09
60670000
32c40794
f88cb33c
4047a026
a00602b4
32dc0007
205c003c
40770a81
d4dc4007
7f5c003b
37c30021
42f24517
23c36026
31c42264
f88c133c
313c44d2
4383fff0
37c4e097
23837f32
0016723c
36c4e0f7
f88c833c
788375c3
e9d227c3
408d5806
60ad6586
456640cd
408640ed
0b0d343c
633c33c4
a5c3f88c
4ac3a683
1d548007
98066100
323c8c8d
23c30010
61002364
8c8d8606
0010323c
236423c3
98066100
323c8c8d
23c30010
61002364
8c8d85e6
0010323c
236423c3
d33c39c4
c5c3f88c
4cc3cd83
1f548007
6100cfd2
8c8d8006
0010323c
236423c3
93e66100
323c8c8d
23c30010
cfd22364
80066100
323c8c8d
23c30010
61002364
8c8d93c6
0010323c
236423c3
60073ac3
61001d54
8c8d8006
0010323c
236423c3
93a66100
323c8c8d
23c30010
61002364
8c8d8006
0010323c
236423c3
93866100
323c8c8d
23c30010
e0072364
2fd21f54
98066100
323c8c8d
23c30010
61002364
8c8d85c6
0010323c
236423c3
61002fd2
8c8d9806
0010323c
236423c3
85a66100
323c8c8d
23c30010
9f5c2364
45c30064
80074983
2fd23054
b8066100
323cac8d
23c30010
61002364
ac8da646
0010323c
236423c3
10542007
b8066100
323cac8d
23c30010
61002364
ac8da626
0010323c
236423c3
8fd20053
b8066100
323cac8d
23c30010
61002364
ac8da4e6
0010323c
236423c3
6100efd2
ac8db806
0010323c
236423c3
a4666100
323cac8d
23c30010
80072364
2fd21054
b8066100
323cac8d
23c30010
61002364
ac8da526
0010323c
236423c3
1054e007
61002fd2
ac8db806
0010323c
236423c3
a4a66100
323cac8d
23c30010
8fd22364
b8066100
323cac8d
23c30010
61002364
ac8da506
0010323c
236423c3
6100efd2
ac8db806
0010323c
236423c3
a4866100
323cac8d
23c30010
80072364
2fd21054
98066100
323c8c8d
23c30010
61002364
ac8da546
0010323c
236423c3
1054e007
61002fd2
8c8d9806
0010323c
236423c3
a4c66100
323cac8d
23c30010
5bc32364
48834bc3
80078037
b0c33b54
7806b284
708d4bc3
0010323c
236423c3
b284b0c3
3bc38146
323c8c8d
23c30010
20072364
b0c31354
7806b284
708d4bc3
0010323c
236423c3
b284b0c3
3bc380a6
323c8c8d
23c30010
b0c32364
7806b284
708d4bc3
0010323c
236423c3
b284b0c3
3bc38126
323c8c8d
23c30010
25f22364
a00702d3
02735d54
b284b0c3
4bc37806
323c708d
23c30010
b0c32364
8086b284
8c8d3bc3
0010323c
236423c3
600738c3
001fe2dc
b284b0c3
3bc39806
323c8c8d
23c30010
b0c32364
60e6b284
708d4bc3
0010323c
236423c3
80c33d53
98068284
8c8d38c3
0010323c
236423c3
828480c3
48c36046
323c708d
23c30010
80172364
1e548007
98066100
323c8c8d
23c30010
61002364
8c8d8106
0010323c
236423c3
61002fd2
8c8d9806
0010323c
236423c3
80666100
323c8c8d
23c30010
85c32364
48c38683
61008fd2
8c8d9806
0010323c
236423c3
82866100
323c8c8d
23c30010
45c32364
80374983
15548007
13542007
b284b0c3
4bc37806
323c708d
23c30010
b0c32364
81e6b284
8c8d3bc3
0010323c
236423c3
600738c3
b0c31354
9806b284
8c8d3bc3
0010323c
236423c3
b284b0c3
4bc36266
323c708d
23c30010
80172364
16548007
16542007
b284b0c3
4bc37806
323c708d
23c30010
b0c32364
81c6b284
8c8d3bc3
0010323c
236423c3
a0070073
c0072954
001642dc
b284b0c3
4bc37806
323c708d
23c30010
b0c32364
8226b284
8c8d3bc3
0010323c
236423c3
90c32a13
78069284
708d49c3
0010323c
236423c3
928490c3
39c38186
323c8c8d
23c30010
38c32364
13546007
928490c3
39c39806
323c8c8d
23c30010
90c32364
62469284
708d49c3
0010323c
236423c3
80078017
2fd21054
38066100
323c2c8d
23c30010
61002364
8c8d81a6
0010323c
236423c3
2954e007
f8066100
323cec8d
23c30010
61002364
2c8d3586
0010323c
236423c3
ec8d6100
0010323c
236423c3
95c66100
323c8c8d
23c30010
61002364
323cec8d
23c30010
61002364
ec8df5e6
0010323c
236423c3
20071ac3
61001c54
8c8d9806
0010323c
236423c3
f4066100
323cec8d
23c30010
61002364
323c8c8d
23c30010
61002364
2c8d3426
0010323c
236423c3
60073cc3
cfd21f54
80066100
323c8c8d
23c30010
61002364
ec8ded66
0010323c
236423c3
6100cfd2
2c8d2006
0010323c
236423c3
8ce66100
323c8c8d
23c30010
15c32364
20071d83
cfd23254
a0066100
323cac8d
23c30010
61002364
ec8de726
0010323c
236423c3
1054c007
20066100
323c2c8d
23c30010
61002364
8c8d8666
0010323c
236423c3
20070073
cfd21054
a0066100
323cac8d
23c30010
61002364
ec8de2c6
0010323c
236423c3
20071ac3
61001c54
8c8d8006
0010323c
236423c3
a7a66100
323cac8d
23c30010
61002364
323c8c8d
23c30010
61002364
ec8de786
0010323c
236423c3
200718c3
61001d54
8c8d8006
0010323c
236423c3
a6a66100
323cac8d
23c30010
61002364
323c8c8d
23c30010
61002364
ec8de5e6
0010323c
236423c3
c0070073
61002b54
2c8d2006
0010323c
236423c3
80a66100
323c8c8d
23c30010
c0072364
61001b54
323c2c8d
23c30010
61002364
ac8da086
0010323c
236423c3
2c8d6100
0010323c
236423c3
e1466100
323cec8d
23c30010
400e2364
40d72097
b8bc6006
02330b3f
600738c3
ffe272dc
24dc2007
c453ffe1
800749c3
ffec12dc
c4dc2007
d793ffea
fc760496
08040f56
50c37016
000761c3
305c2154
6ed20824
10f8301c
0000311c
8c4c6c0c
40a6000c
66f0301c
0017311c
055c4664
0ed20864
10f8301c
0000311c
8c4c6c0c
454616c3
66f0301c
0017311c
0e564664
00000804
10fc301c
0000311c
6c6c6c0c
36640006
00000804
ff961016
226440c3
00074037
400d1254
1561235c
235c402d
404d1569
1e24335c
4000341c
01c366f2
0030143c
0b3f08bc
08560196
00000804
2f5c30c3
233c0021
01c300df
f4bc13c3
08040b3e
fd967016
51c360c3
226443c3
208540b7
24bc42c6
3f5c0b44
3f5c0041
80770005
0050063c
400615c3
40bc35c3
03960b44
08040e56
0136f016
70c3fd96
82c351c3
829763c3
01213f5c
208560b7
34c342c6
0b4424bc
00413f5c
00053f5c
073c8077
16c30050
35c328c3
0b4440bc
80760396
08040f56
50c3f016
62c371c3
6eac600c
26546007
8eac740c
17c305c3
748c26c3
00074664
1f871e15
1f87f654
1f4706d4
1f671754
01f31694
06541fc7
07741fc7
0f941fe7
001c01b3
0173febd
1e24355c
00936f72
1e24355c
355c7072
1fe61e27
08040f56
40c33016
10f8301c
0000311c
205c6c0c
ac4c0444
04c9305c
312c09a0
301c4186
311c6688
56640017
0800343c
0447345c
345c60a6
600604a7
04c5345c
04cd345c
08040c56
50c37016
6ecc600c
35946007
740c0873
0444255c
05c38ecc
0484355c
26c32980
466474ac
15150007
25541f87
04d41f87
30941f67
1fa70113
201c0654
1fc7feb9
05532994
1e24355c
355c6f72
04531e27
0464255c
03e432c3
201c04f4
0393fe7d
0484355c
355c6c00
355c0487
6c200464
0467355c
0464655c
ca94c007
0487655c
04c1355c
68d223c3
b4bc05c3
26c30b44
201c0073
02c3fecc
08040e56
51c37016
280c43c3
0040313c
001c680f
4157ff7c
36e462c3
74800ab4
009f233c
03c3500d
30bc2117
00060b3f
08040e56
02641016
031c1264
319400cc
00a9131c
000d52dc
00a9131c
228711b4
000cf2dc
05b42287
24dc2267
1673000e
165422a7
00a8131c
000db4dc
131c1593
32dc00ab
131c000d
0a1400ab
00ac131c
000c92dc
00ad131c
000cb4dc
45f20073
408737f3
001bd2dc
24dc4027
3713000c
00c0031c
000bd4dc
45b42507
71dc24e7
21a70009
0008b2dc
27b421a7
72dc20c7
20c7000a
206711b4
000992dc
05b42067
04dc2047
1253001a
02dc2087
20a70009
001994dc
21271173
000832dc
07b42127
7e5420e7
e4dc2107
0f530018
78542147
84dc2187
0c530018
5d542267
0bb42267
5c5421e7
5a1421e7
55542227
a4dc2247
0a330017
67b42487
71342467
24dc2287
09330017
6e542747
1fb42747
5e5425c7
0bb425c7
54542567
4f142567
5f542587
04dc25a7
06930016
38542627
07b42627
315425e7
64dc2607
05b30015
2e542647
04dc26e7
0a330015
00a7131c
131c10b4
3f3400a6
00a0131c
001450dc
00a1131c
131c2035
e0dc00a4
07930013
00ac131c
131c2754
06b400ac
00a9131c
001335dc
313c0633
6027f520
0012d5dc
40670333
24d32f94
2c944007
40672473
24130b94
e2dc4007
40c70011
23532394
82dc4007
40c70011
22931d94
089440c7
40472233
21d31794
c2dc4047
40670010
21131194
62dc4087
40270010
20530b94
08944047
40871ff3
1f930594
a2dc4087
031c000f
82dc00c0
031c000f
42dc00cc
131c000f
61b4009d
009c131c
000d51dc
92dc2727
2727000c
22c72cb4
000d82dc
14b422c7
82dc20a7
20a7000c
204708b4
000c32dc
84dc2087
17d3000d
c2dc20e7
2147000b
000d14dc
266716f3
000a62dc
08b42667
22dc2587
25e70009
000c54dc
26871573
000ba2dc
e4dc26a7
1493000b
72dc2ce7
2ce70008
27a714b4
0009d2dc
08b427a7
82dc2767
27870009
000ad4dc
28271273
000912dc
64dc28a7
11f3000a
0088131c
0008c2dc
0088131c
2d6708b4
131c6e54
84dc0084
0fd30009
f740313c
25dc6027
0b530009
00be131c
131c7854
1cb400be
00ab131c
131c0bb4
4c3400aa
009f131c
131c6635
7e1400a8
131c08f3
08b400b5
00b2131c
131c3f34
741400ae
131c07b3
709400ba
131c0af3
2c5400e8
00e8131c
131c15b4
265400e5
00e5131c
131c08b4
485400c0
00c4131c
08f35d94
00e6131c
131c1954
569400e7
131c02b3
3a5400fa
00fa131c
131c05b4
4c1400f8
131c0673
305400fc
00fc131c
131c2d14
429400fd
323c0533
333c0056
7fe50b0d
f88c033c
40270753
323c3554
fed30046
30544007
40270006
05533094
2a544007
40270006
04932a94
24544007
40270006
03d32494
1e544007
40270006
03131e94
10944007
323c02f3
fb530b0d
12544007
105440c7
40270006
01531094
40c74bd2
323c0954
f9530016
40270006
02c30694
00260093
00060053
08040856
0336f016
40c3fc96
72540007
70544007
6ef42007
5dc4601c
0017611c
70093810
59c36037
15a273c3
341c30c3
63d20001
e037e405
00010f5c
00070064
80255254
35940547
20073fe5
200704d4
03931554
009f343c
780c6077
eea2a057
341c37c3
63d20001
a077a405
00213f5c
65473064
03c3ea54
01c30133
30e400f3
65c72754
40253754
b80c0053
60b76809
87c3f5a2
0001841c
65d238c3
37c3e097
60b76405
00413f5c
60073064
0213e994
a0f7a809
eea2780c
341c37c3
63d20001
a0f7a405
00613f5c
03e43064
68081394
0b0d333c
7f3233c4
20074980
3fe504f4
a0942007
303c0809
7fe50b0d
03c37f32
00060053
c0760496
08040f56
21c3ff96
41872264
000862dc
11b44187
3d544047
06b44047
24544007
1f944027
40870533
40874754
41673914
09331894
f2dc4207
4207000b
41c70ab4
000812dc
1544105c
a5dc41c7
0e73000a
4e5442c7
02dc46e7
4287000d
000bb2dc
fe76001c
305c1fb3
233c1544
60720014
1e544007
305c1dd3
133c1544
20070024
000e84dc
085b323c
1547305c
1d1301c3
1544305c
0044233c
4ad26272
305c1b53
233c1544
40070084
000d44dc
305c6372
02c31547
305c1ab3
233c1544
64720104
18f357d2
1544205c
0204323c
14dc6007
4572000c
1547205c
1e24305c
0010341c
323c64d2
0e730044
0024323c
205c0e13
323c1544
60070404
000ac4dc
205c4672
323c1547
60070204
000a72dc
0804323c
52dc6007
1413000a
1544205c
0804323c
74dc6007
32c30009
305c6772
341c1547
09b30004
1004213c
687231c3
b8544007
205c1113
323c1544
60072004
000824dc
205c4972
323c1547
60070204
305c1294
13c315d9
20373f85
00013f5c
09356047
1e24305c
111c2006
31834000
6c546007
0804323c
6b946007
15f9305c
67546027
15d9005c
63540027
5e9400e7
313c0c13
60074004
31c35694
305c6a72
341c1547
01b30020
1544205c
8004323c
49946007
6b7232c3
1547305c
0002341c
47946007
205c0873
32c31544
1000341c
39946007
6c7232c3
1547305c
2000341c
fe77001c
35946007
205c06b3
32c31544
2000341c
27946007
1e24305c
4000341c
32c365f2
305c6d72
105c1547
313c1e24
213c0104
67d24004
305c4cf2
341c1544
00d30200
305c46f2
341c1544
6ed20800
341c31c3
6dd24000
1544305c
305c6d72
00f31547
fe75001c
001c00b3
0053fe8b
01960006
00000804
28d220c3
1d84005c
0010303c
1d87325c
005c00f3
303c1da4
325c0010
08041da7
60e6fe96
1d39105c
402521c3
1f5c4037
20770001
00212f5c
1d3d205c
7fe525f2
7fe71fe5
0296f094
00000804
41c31016
15e9205c
15c9305c
12946027
15a3105c
3410341d
18946007
21e44025
21c30234
1e24305c
2000341c
48806cd2
60470153
205c0894
305c15b3
614715c1
41050254
42e40006
001c0334
0856fe89
00000804
50c37016
21c342c3
20062264
00d301c3
d4a232c3
03a33603
14e42025
0e56fa74
00000804
303c3016
8d20fd60
fd50303c
ad206ca0
f90c343c
003f341c
233c6e00
353c310c
341cf90c
6e80003f
49a06652
343c0006
62d203f4
08000026
353c2006
62d203f4
00a02026
08040c56
40c3f016
62c351c3
e15703c3
323c480c
37e40020
352229b4
0010323c
55a2780f
780f6025
1387245c
145c51c3
400f13a7
06942047
1e24345c
345c7072
600c1e27
345c66f2
71721e24
1e27345c
200604c3
0b3eeabc
780c0bd2
1de4145c
07e40c80
180f03b4
501c0073
05c3ff7c
08040f56
08040006
5dc8001c
0017011c
00000804
63e0001c
0017011c
00000804
080406c6
ff967016
602c52c3
15e1205c
0a95235c
c046602c
0a8d635c
03d38026
305c4429
23e415e1
44091794
40474037
c0171754
408726c3
40170954
60a732c3
40170554
60c732c3
602c0794
00016f5c
0a8d635c
804500b3
45e42045
0196e214
08040e56
005c30c3
135c1e59
40861e61
0b453cbc
0b0d303c
033c7fe5
0804f88c
0336f016
80c3ff96
52c391c3
c80c73c3
a2dc6007
67220009
00163f5c
0010163c
2f5c280f
323c0013
37e40010
0008d5dc
940f8500
0b3ed2bc
20540007
60457320
25dc37e4
19c30008
1f3c0600
3ebc0020
740c0b3f
0020133c
2f5c340f
67200013
37e46d00
08c371b4
2c8039c3
0b49a8bc
4f5c740c
6e000013
540c740f
0020323c
37e46f20
19c361b4
1f3c0500
3ebc0020
740c0b3f
740f6045
2f5c6f20
6d000013
203537e4
540c0a33
0020323c
37e46f20
39c34bb4
1fc30d00
0b3f3ebc
233c740c
540f0020
00031f5c
6c806b20
3cb437e4
740f6880
00132f5c
7fc532c3
3f5c6ca0
3f5c0016
60070013
48c3df94
0744345c
10546007
6ed26c0c
0764345c
6c0c6bd2
345c69d2
40261e24
101b323c
1e27345c
08c301b3
0b3ec4bc
08c309d2
1e24305c
323c4046
305c101b
08c31e27
eabc2006
30c30b3e
740c6bd2
115c18c3
6c801de4
0006740f
001c0073
0196feb8
0f56c076
00000804
00d1301c
1a5402a7
0ad402a7
00b8301c
14540207
0208301c
0e940267
301c01f3
030700d2
301c0b54
032700d3
301c0754
02e7020e
301c0354
03c3fea1
00000804
0007ff96
004c2754
24540007
6306016c
031c6037
205400d2
00d2031c
62060cb4
031c6037
185400b8
603762a6
00d1031c
02531194
60376266
0208031c
62e60d54
031c6037
0854020e
60376326
00d3031c
60060354
3f5c6037
03c30001
08040196
fd96f016
236421c3
1e24505c
2007202c
000852dc
600675c3
0400311c
65007383
20772c89
60b76ca9
400665c3
0080211c
80066283
46c3c4f2
8026e2f2
00213f5c
2f5c03c3
12c30041
3cbc4006
03d20b45
64548007
00213f5c
2f5c03c3
12c30041
3cbc4026
08d20b45
200635c3
0040111c
60073183
2f5c5354
02c30021
00413f5c
404613c3
0b453cbc
35c308d2
111c2006
31830020
42546007
00212f5c
3f5c02c3
13c30041
3cbc4066
03d20b45
3654e007
00211f5c
2f5c01c3
12c30041
3cbc4086
00070b45
3f5c2b94
03c30021
00412f5c
40a612c3
0b453cbc
c00703d2
3f5c1f54
03c30021
00412f5c
40c612c3
0b453cbc
00076026
60061454
111c2206
51830200
211c4006
12c30200
029451e4
133c6026
20370016
00013f5c
60060053
039603c3
08040f56
f996f016
61c370c3
323c42c3
331cf820
42b40082
0200063c
01a01f3c
0b3f3ebc
00d30f5c
fbe0343c
03e43364
2f3c35b4
023c01c0
3c0cfc7e
6006b800
363c6037
60770220
40f700b7
0484215c
415c4137
07c30464
263c16c3
353c0100
46640220
000750c3
41571e74
00d33f5c
17d423e4
15f44767
004703d2
463c1494
7c4c0220
2710033c
0260163c
b0bc4606
538b08cb
0a76275c
501c00d3
0073fe71
fe72501c
079605c3
08040f56
50c3f016
63c342c3
305ce157
341c1e24
6ff24000
480c06c3
40a62500
08cbb0bc
60a5700c
063c700f
17c30030
0b3f3ebc
233c780c
355c820b
23e41563
255c1b54
323c1e24
65f20104
1e99355c
12356027
2104323c
0210331c
355c0594
60671e91
32c30935
4000341c
22546007
62c77809
3c0b1f94
47a3255c
1118301c
0000311c
6c4c6c0c
023523e4
323c23c3
001c0660
13e4feab
18090fd4
7d8530c3
fec9001c
08b46067
255c4006
00061e0d
001c0073
0f56feba
00000804
0136f016
80c3ff96
42c351c3
c80c73c3
28356047
00200f3c
40462700
08cbb0bc
233c700c
500f0020
00113f5c
00fe331c
3f5c1c94
331c0019
045400ff
00fd331c
35221494
500f4025
6b2027d2
37e46c80
650009b4
4026700f
215c18c3
00061e6d
001c00d3
0073feb8
feba001c
80760196
08040f56
0136f016
50c3fd96
62c381c3
880c73c3
fe7a001c
4801155c
92dc2007
6067000b
000b49dc
0e0038c3
00401f3c
0b3f48bc
233c780c
580f0040
60456a20
55dc37e4
38c3000a
1f3c0d00
3ebc00a0
780c0b3f
780f6045
00532f5c
6d006e20
55dc37e4
355c0009
231c1371
33350100
10546007
10f8301c
0000311c
8c4c6c0c
0b44055c
4726352c
65f4301c
0017311c
301c4664
311c10f8
6c0c0000
0f5c8c0c
352c0053
301c4726
311c65f4
46640017
055c0037
0bf20b47
16e0353c
0b47355c
00013f5c
1375355c
0c731066
455c8026
03331375
10546007
10f8301c
0000311c
8c4c6c0c
0b44055c
4726352c
65f4301c
0017311c
20064664
1375155c
16e0353c
0b47355c
00532f5c
30544007
0b44055c
980c38c3
b0bc2e00
3f5c08cb
580c0053
580f4980
0b66355c
155c2057
455c14a7
89d247c4
155c05c3
255c0b44
355c0b63
466447e4
1e24355c
355c6b72
544c1e27
00533f5c
3c0513c3
0b44355c
0500023c
44062c80
08cbb0bc
255c0073
05c30b66
eabc2006
06d20b3e
455c780c
6e001de4
2006780f
4805155c
00730006
feb8001c
80760396
08040f56
0336f016
50c3fe96
305c91c3
341c1e24
e1a64000
e0a662f2
163cc086
2077080c
00216f5c
fa1467e4
10f8301c
0000311c
09c36c0c
0464155c
8c0c4080
352c0b00
301c4186
311c6650
46640017
106620c3
34544007
82c37ba0
255c8384
46d20464
155c08c3
b0bc0444
155c08cb
200704c1
301c1354
311c10f8
6c0c0000
0444255c
355c8c4c
09a004c9
4186352c
6650301c
0017311c
00264664
04c5055c
e037fba0
00011f5c
04cd155c
0447855c
055c29c3
68000464
04a7355c
02960006
0f56c076
00000804
201c3016
2007ff53
305c0e74
205c04a4
6d200464
063431e4
0b4d26bc
00075066
40060274
0c5602c3
00000804
0136f016
50c3fe96
305c72c3
341c1e24
42064000
62f24077
e0076077
20070374
001c0415
09d3ff53
818487c3
10f8301c
0000311c
8c0c6c0c
02c34057
352c0884
301c41a6
311c6664
46640017
106660c3
3854c007
63d26057
d9807e65
776ce8d2
57ac06c3
27c32d00
08cbb0bc
03e1355c
12546007
10f8301c
0000311c
576c6c0c
355c8c4c
09a003e9
41a6352c
6664301c
0017311c
40264664
03e5255c
68d26057
60377e65
00013f5c
03ed355c
2f5c00b3
255c0021
d76f03ed
600617d1
f78f77af
029603c3
0f568076
00000804
50c3f016
638c71c3
8d2043ac
6e2063cc
38748007
36746007
c007c620
63e433f4
24c308f4
0b4d9ebc
106630c3
2c746007
57ac89d2
776c47d2
2d0003c3
b0bc24c3
600608cb
978f77af
05c3776c
2d00578c
84bc26c3
1fe70b44
001c0494
0293fecc
febd031c
06e41154
001c04f4
0193fe88
6100578c
37e4778f
00060314
d82000b3
001cfc93
0f56feb8
00000804
50c37016
638c43ac
313ccd20
7fe50b0d
63d27f32
29d4c0a7
c0076ad2
776c08f4
0640053c
26c32d00
08cbb0bc
10f8301c
0000311c
576c6c0c
155c8c4c
08a003e9
41a6352c
6674301c
0017311c
353c4664
776f0640
77cf60a6
155c2006
155c03e5
600603ed
d78f77af
08040e56
40c31016
1a540007
0040303c
6006600f
0827305c
010c021c
4b862006
0891b0bc
1680043c
44062006
0891b0bc
16c0343c
0be7345c
345c6006
08560c47
00000804
ff961016
203740c3
2587205c
20060085
0b4e80bc
1900043c
80bc2006
60060b4e
345c700f
345c24c7
345c2467
345c2527
345c2547
3f5c2567
345c0001
600625a5
25ad345c
345c6006
345c2507
345c25c7
345c25f5
345c25fd
345c2605
345c260d
345c2615
345c261d
60062625
2647345c
2667345c
2685345c
268d345c
345c6006
345c26a7
345c26c7
345c26e5
600626ed
25e6345c
08560196
00000804
0736f016
50c3e296
0b44605c
0180af3c
20060ac3
b0bc4786
155c0891
1f5c1561
255c00c5
2f5c1569
355c00cd
3f5c1e59
155c00d5
1f5c1e61
744c00dd
01c00f3c
2710133c
b0bc4606
1abc08cb
1f3c0b44
16bc04c0
355c0b3f
333c1e44
3f5c0acb
763c0286
07c30220
47861ac3
08cbb0bc
07803f3c
00be201c
fe7e233c
963c540c
863c0100
20260e00
e0772037
20b72786
325c60f7
61370484
0464425c
16c305c3
38c329c3
01774664
48940007
78856757
0082331c
301c0535
6177fe72
07c307f3
47861ac3
08cbeabc
35540007
05404f3c
2f5c04c3
12c300a1
b0bc4406
06c30891
420614c3
08cbeabc
25540007
14c309c3
eabc4206
000708cb
08c31e54
440614c3
08cbeabc
17540007
03a30f5c
0200163c
0b3f08bc
323c4757
355c0420
231c0b66
0cd400bd
033c7900
18c30220
b0bc4406
009308cb
fe70201c
01574177
e0761e96
08040f56
305c10c3
600748c4
02331094
033c644c
121c0500
440600fc
08cbeabc
0b0d303c
033c7fe5
01b3f88c
01730026
0b63305c
305c7cf2
341c1e24
03c30800
e7946007
00000804
0136f016
01c340c3
13c362c3
1e24345c
1000341c
62f2a186
201ca486
51e4feb8
380c3d94
1de4745c
6e806780
ff7c201c
87c3e197
32b438e4
4af241d7
306c0080
eabc25c3
201c08cb
0007fed0
f80c2794
245c7780
6d001de4
345c780f
233c1e24
033c0104
4ed24004
345c60c6
00071e6d
e1461494
1e7d745c
245c4026
20c31e85
612601b3
1e75345c
e14608d2
1e7d745c
345c6026
00531e85
02c34006
0f568076
00000804
40c37016
a58060a5
ffb0623c
033c606c
15c31680
dabc26c3
706c0b1d
1c80033c
26c315c3
0b05a6bc
d2bc04c3
30c30b3e
19546007
033c706c
15c32240
aabc26c3
00070b1d
706c1094
2900033c
26c315c3
0b1d4abc
706c08f2
35c0033c
26c315c3
0b1d7abc
08040e56
0136f016
305c50c3
341c1e44
66d20100
0b4eeebc
000760c3
355c3f94
833c0b63
733c0060
05c300f0
88bc17c3
60c30b4d
32940007
0444355c
0464255c
04c38d00
408618c3
4abc35c3
740c0b44
04a4035c
0090143c
0b3f16bc
0b63055c
00d0143c
0b3f08bc
00f0043c
0b44155c
0b63255c
08cbb0bc
14c305c3
36c327c3
0b5004bc
0af260c3
0464355c
355c6f80
05c30467
0b44d6bc
06c360c3
0f568076
00000804
60c37016
88bc2126
50c30b4d
20940007
0444365c
0464265c
04c38d00
41c615c3
4abc36c3
06c30b44
412614c3
04bc35c3
50c30b50
60a60df2
1e6d365c
0464365c
365c6125
06c30467
0b44d6bc
05c350c3
08040e56
40c3f016
0b3ed2bc
05d2c086
4c2b702c
c0c562c3
1e24345c
211c4006
32836000
60070006
763c5494
04c30090
88bc17c3
00070b4d
345c4c94
245c0444
ad000464
16c305c3
34c341a6
0b444abc
752d6026
1e59345c
00c0331c
345c0894
606715e1
68060494
0073754d
554d4026
d2bc04c3
61660b3e
13540007
0c2b702c
00b0153c
0b3f08bc
053c702c
133c00d0
4c2b1300
08cbb0bc
4c2b702c
61a532c3
35800006
0b3f08bc
15c304c3
600627c3
0b5004bc
345c0ef2
6f800464
0467345c
1e44345c
0008341c
04c364f2
0b44d6bc
08040f56
40c37016
62c351c3
033c606c
dabc1680
706c0b1d
1c80033c
26c315c3
0b05a6bc
d2bc04c3
30c30b3e
19546007
033c706c
15c32240
aabc26c3
00070b1d
706c1094
2900033c
26c315c3
0b1d4abc
706c08f2
35c0033c
26c315c3
0b1d7abc
08040e56
40c37016
ffc0513c
0040623c
033c606c
15c31680
dabc26c3
706c0b1d
1c80033c
26c315c3
0b05a6bc
d2bc04c3
30c30b3e
19546007
033c706c
15c32240
aabc26c3
00070b1d
706c1094
2900033c
26c315c3
0b1d4abc
706c08f2
35c0033c
26c315c3
0b1d7abc
08040e56
50c37016
0564005c
13540007
10f8301c
0000311c
8c4c6c0c
44c6352c
6308301c
0017311c
60064664
0567355c
0587355c
05a4055c
13540007
10f8301c
0000311c
8c4c6c0c
44c6352c
6308301c
0017311c
60064664
05a7355c
05c7355c
0007158c
d5ac1d54
0454c147
1594c4a7
e6bc0093
00730b1c
0ad2b6bc
10f8301c
0000311c
8c4c6c0c
352c158c
301c26c3
311c6308
46640017
75af6006
0e56758f
00000804
fe96f016
26bc50c3
03640b96
0460703c
1e44355c
0200341c
40774406
744c6ed2
0381335c
001c6077
6407feb8
000915dc
32c34057
fd807c05
101c05c3
88bc0080
00070b4d
000854dc
0444355c
0464255c
06c3cd00
404617c3
4abc35c3
355c0b44
792d1561
1569255c
355c594d
341c1e24
463c0400
600700b0
14cc1b94
605714c3
442523c3
0b1bf6bc
62940007
033c744c
14c30300
b0bc4406
2f5c08cb
265c0021
744c015d
0500033c
02c0163c
744c0233
133c04c3
44060300
08cbb0bc
00213f5c
015d365c
063c744c
133c02c0
40570500
08cbb0bc
32c34057
255c6585
59a11e59
32c34057
255c65a5
59a11e61
13c36057
255c25c5
60061e24
0008311c
40372383
23c36057
601745e5
7ba663d2
3f5c0073
78a10001
0090473c
390005c3
0b9600bc
0464355c
355c6e00
05c30467
24c316c3
04bc6006
0cf20b50
255c4046
355c1e6d
341c1e44
64f20008
d6bc05c3
02960b44
08040f56
0136f016
80c3e996
62c371c3
eebc0fc3
a0060b00
0fc300f3
26c317c3
0b05a6bc
58e4a025
1796f974
0f568076
00000804
0736f016
40c3fc96
801ca1c3
811c10f8
28c30000
901c680c
911c6390
ac0c0017
20060b86
39c344c6
70c35664
680c28c3
0b86ac0c
44c62006
566439c3
706c50c3
133c07c3
4b861c80
08cbe6bc
504c706c
1c80033c
2710123c
a6bc4606
706c0b05
1c80033c
6330101c
0017111c
a6bc4606
706c0b05
1c80033c
66bc1fc3
706c0b25
1c80033c
0abc17c3
05c30b24
0b00eebc
05c3704c
2710133c
a6bc4606
05c30b05
6360101c
0017111c
a6bc4606
05c30b05
42061fc3
0b05a6bc
1ac305c3
0b055cbc
680c28c3
07c38c4c
44c62006
466439c3
680c28c3
05c38c4c
44c62006
466439c3
e0760496
08040f56
0736f016
40c3fc96
62c3a1c3
10f8701c
0000711c
901c7c0c
911c65b8
ac0c0017
20060b86
39c344c6
80c35664
ac0c7c0c
20060b86
39c344c6
50c35664
08c3706c
1c80133c
e6bc4b86
706c08cb
1c80033c
408616c3
0b05a6bc
504c706c
1c80033c
2710123c
a6bc4606
706c0b05
1c80033c
6330101c
0017111c
a6bc4606
706c0b05
1c80033c
66bc1fc3
706c0b25
1c80033c
0abc18c3
05c30b24
0b00eebc
05c3704c
2710133c
a6bc4606
05c30b05
6360101c
0017111c
a6bc4606
05c30b05
42061fc3
0b05a6bc
1ac305c3
0b055cbc
8c4c7c0c
200608c3
39c344c6
7c0c4664
05c38c4c
44c62006
466439c3
e0760496
08040f56
0136f016
80c3e896
62c371c3
ecbc0fc3
a0060b1d
0fc300f3
26c317c3
0b1ddabc
58e4a025
1896f974
0f568076
00000804
0736f016
40c3fb96
801ca1c3
811c10f8
28c30000
901c680c
911c63a4
ac0c0017
20060c06
39c344c6
70c35664
680c28c3
0c06ac0c
44c62006
566439c3
706c50c3
133c07c3
4c061680
08cbe6bc
504c706c
1680033c
2710123c
dabc4606
706c0b1d
1680033c
6330101c
0017111c
dabc4506
706c0b1d
1680033c
4ebc1fc3
706c0b25
1680033c
0ebc17c3
05c30b24
0b1decbc
05c3704c
2710133c
dabc4606
05c30b1d
6360101c
0017111c
dabc4506
05c30b1d
42861fc3
0b1ddabc
1ac305c3
0b1dcabc
680c28c3
07c38c4c
44c62006
466439c3
680c28c3
05c38c4c
44c62006
466439c3
e0760596
08040f56
9a96f016
61c340c3
0f3ca06c
153c0cc0
201c2900
e6bc00cc
0fc308cb
35c0153c
00cc201c
08cbe6bc
1e24345c
1000341c
0100763c
2c546007
1c80053c
66bc16c3
706c0b25
1680033c
4ebc17c3
04c30b25
0b3ed2bc
24540007
033c706c
163c2240
00bc0240
00070b25
706c3394
2900033c
0440163c
0b1d3abc
2a940007
033c706c
163c35c0
6abc0740
0ad20b1d
04c30433
90bc16c3
04c30b52
94bc17c3
04c30b53
0b3ed2bc
600730c3
706c1354
2900033c
0cc01f3c
00cc201c
08cbe6bc
033c706c
1fc335c0
00cc201c
08cbe6bc
66960006
08040f56
0736f016
40c3fb96
62c3a1c3
10f8701c
0000711c
901c7c0c
911c65c4
ac0c0017
20060c06
39c344c6
80c35664
ac0c7c0c
20060c06
39c344c6
50c35664
08c3706c
1680133c
e6bc4c06
706c08cb
1680033c
408616c3
0b1ddabc
504c706c
1680033c
2710123c
dabc4606
706c0b1d
1680033c
6330101c
0017111c
dabc4506
706c0b1d
1680033c
4ebc1fc3
706c0b25
1680033c
0ebc18c3
05c30b24
0b1decbc
05c3704c
2710133c
dabc4606
05c30b1d
6360101c
0017111c
dabc4506
05c30b1d
42861fc3
0b1ddabc
1a3c05c3
cabc0100
7c0c0b1d
08c38c4c
44c62006
466439c3
8c4c7c0c
200605c3
39c344c6
05964664
0f56e076
00000804
50c33016
204c31c3
6cd22dd2
00fc021c
44062a05
08cbb0bc
235c744c
255c0381
144c08e5
17540007
10f8301c
0000311c
8c4c6c0c
352c000c
301c4426
311c66d0
46640017
4006744c
144c4c0f
02a4101c
0b06b8bc
10f8301c
0000311c
8c4c6c0c
352c144c
301c4426
311c66d0
46640017
744f6006
08040c56
0336f016
71c340c3
5d540007
5df0101c
0017111c
089298bc
601c06d2
611c5df0
03730017
101c04c3
111c5df8
98bc0017
06d20892
5df8601c
0017611c
04c301d3
5dfc101c
0017111c
089298bc
05d260c3
5dfc601c
0017611c
901ca006
911c64b8
801c0017
811c63e0
29c30017
37e46a81
38c32694
80078e81
c0072254
04c31b94
5df0101c
0017111c
089298bc
17940007
101c04c3
111c5df8
98bc0017
0ff20892
101c04c3
111c5dfc
98bc0017
07f20892
04c30193
98bc16c3
07f20892
531ca085
d49400d8
00530006
c07604c3
08040f56
61c37016
000750c3
a12c1254
942c0213
0ebc04c3
30c30892
04c33364
26c313c3
0b472ebc
002603d2
b40c0093
05c3b1f2
08040e56
41c31016
0b499abc
04c330c3
4a0613c3
0892e6bc
08040856
3f36f016
70c3f296
a6bc41c3
d0c30b49
83f2e2d2
1933a006
300964c3
42dc2007
04c3000c
5e00101c
0017111c
2abc4066
01640892
82dc0007
a006000b
b5c395c3
c5c3a5c3
101c06c3
111c5e04
98bc0017
80c30892
06c307f2
08920ebc
136410c3
28c30073
06262b20
0b3ebebc
0f3c40c3
16c30070
e6bc24c3
86270892
86060294
00703f3c
2e212006
63c38006
06c30ef3
63e0201c
0017211c
4a1d123c
3ebc4626
00070bfe
06c36a94
5df0101c
0017111c
089298bc
00cc101c
00072037
06c32194
5e08101c
0017111c
089298bc
00d0301c
00076037
06c31594
5df8101c
0017111c
089298bc
06c30af2
5dfc101c
0017111c
089298bc
04d20037
00c0201c
19c34037
2f5c7c80
4c8d0001
0010293c
101c7d00
111c64b8
113c0017
2c8d489d
0010923c
4ef22ac3
00700f3c
5e0c101c
0017111c
089298bc
a01c05d2
5ac30001
4f3c0473
04c30070
5e14101c
0017111c
089298bc
c01c05d2
5cc30001
3bc302b3
11946007
101c04c3
111c5e18
98bc0017
09f20892
0001b01c
00d35bc3
4de48025
00538974
28c3a026
683c44d2
ebb30010
6026aed2
0a85375c
0006975c
1ac307c3
3cc32bc3
0b3fb8bc
a0260053
0e9605c3
0f56fc76
00000804
40c31016
043c89d2
8cbc03c0
145c0ba0
28bc1e61
08560b55
00000804
0336f016
81c350c3
301c92c3
311c10f8
6c0c0000
001c8c0c
200600cc
301c44c6
311c65a8
46640017
a3d270c3
11940007
10f8301c
0000311c
8c4c6c0c
200607c3
301c44c6
311c65a8
46640017
07b3d066
133c746c
201c2900
e6bc00cc
355c08cb
341c1e24
63c31000
05c367d2
29c318c3
0b9b1abc
355c60c3
341c1e24
6bf21000
18c305c3
04bc29c3
05c30b53
29c318c3
0b5472bc
d2bc05c3
09d20b3e
033c746c
17c32900
00cc201c
08cbe6bc
10f8301c
0000311c
8c4c6c0c
200607c3
301c44c6
311c65a8
46640017
c07606c3
08040f56
0f36f016
70c3f396
a2c391c3
636463c3
0281005c
62dc0007
875c000c
831c15c1
24540007
0007831c
831c09b4
0e540001
0004831c
000b74dc
831c01f3
1c540008
0009831c
000af4dc
1e2c0bd3
9ebc36c3
a0060aa1
301c1533
311c10fc
6c0c0000
1e4c8eac
466436c3
1e6c00b3
68bc36c3
50c30b1e
bf3c1333
0bc301b0
41a62006
0891b0bc
200607c3
0b48dabc
01f01f3c
0b3f16bc
02300f3c
ffb01a3c
b0bc4066
bf0608cb
15b3075c
19807420
02601f3c
0b3f08bc
02804f3c
173c04c3
40863a80
08cbb0bc
02c00f3c
3a00173c
b0bc28c3
275c08cb
3e6c15b3
8037b520
60776186
09c37920
60b76180
bf5c40f7
41a60087
01c34177
0080193c
00802a3c
1ebc7700
08f30b1e
01b08f3c
200608c3
b0bc41a6
07c30891
dabc2006
1f3c0b48
16bc01f0
0f3c0b3f
1a3c0230
4066ffb0
08cbb0bc
075cbf06
742015b3
1f3c1980
08bc0260
4f3c0b3f
04c30280
3a80173c
b0bc4086
0f3c08cb
173c02c0
41063a00
08cbb0bc
15b3275c
b5203e6c
61868037
79206077
618009c3
40f760b7
00878f5c
417741a6
193c01c3
2a3c0080
77000080
0a9e70bc
07c350c3
0b48eabc
218604c3
0b06b8bc
501c0073
05c3fec6
f0760d96
08040f56
3f36f016
50c3f996
d2c381c3
cf5ca3c3
9f5c0244
000702a4
000be2dc
06f209c3
92dc2007
68f2000b
200716d3
000b44dc
14dc6007
b55c000b
3c3c15e9
4bc30050
355cee00
c00615c9
6027c0b7
455c2394
355c15a3
341c1e24
63c32000
11546007
8207fe00
0009b5dc
6af239c3
1f3c14cc
24c300c0
0b1bf6bc
24dc0007
64c30009
0010373c
ffc0273c
2240341d
80b79120
355cf180
604715c9
355c1794
614715c1
c1060254
15b3255c
3ba432c3
ef006f80
600739c3
0f3c6e94
153c00c0
41063a00
08cbb0bc
49c30093
63948007
66b47de4
ffb0373c
936493c3
19c308c3
02613f5c
35c323c3
0b4424bc
cfd280a6
220606c3
0b3ebebc
083c30c3
1f3c0050
23c300c0
08cbb0bc
0050463c
0a0028c3
2cc31ac3
08cbb0bc
03c364d7
0c9402c7
4ad24517
18c305c3
00502c3c
04bc36c3
00070b50
3cc33794
355c3180
602715c9
0bc30e94
40066400
718048c3
00410f5c
40250d21
04c38097
f93520e4
15c9355c
10546047
0050363c
803784d7
c077c006
05c3960c
288028c3
3cc34980
00074664
383c1194
05c30050
23c313c3
06bc39c3
08f20b57
00d307c3
ff53001c
001c0073
0796ff7c
0f56fc76
00000804
0736f016
50c3fa96
1e24305c
4004233c
44d24177
08e1105c
742c2177
fe8d001c
82dc6007
4007000f
255c1a54
40070b63
00061654
0b44155c
6abc752c
10c30b94
72dc0007
201c000e
150008f0
38bc552c
00270b93
000df4dc
21772006
8c0b742c
200605c3
0b93f8bc
44dc0007
343c000d
41570270
05c38d00
0b96acbc
02d20364
943c9000
05c30090
eabc2026
03d20b3e
06f0943c
19c305c3
0b4d88bc
a4dc0007
355c000b
155c0444
cc800464
14c306c3
35c34026
0b444abc
1561255c
355c592d
794d1569
1563155c
1576155c
1e91255c
12944007
00b0463c
14c314cc
f6bc4406
00070b1b
000974dc
033c744c
14c30100
b0bc4406
3f5c08cb
365c00a1
8586015d
2dd22157
02c0063c
0fc0153c
08e1255c
08cbb0bc
08e1255c
858542c3
0c0b742c
08bc3a00
80450b3f
1a00742c
0040133c
b0bc4c0b
742c08cb
70802c0b
59a14026
155c6025
40061e24
0008211c
21371283
0010733c
3ba624d2
009339a1
00812f5c
05c359a1
40bc3b80
40c30b96
05c34364
eabc2026
30c30b3e
39540007
ffb0373c
a01cee00
a11c10f8
1ac30000
8c0c640c
352c07c3
301c44c6
311c63d0
46640017
000780c3
163c3654
27c30050
08cbb0bc
42c6e037
60264077
200660b7
05c320f7
29c316c3
debc38c3
90c30b57
680c2ac3
08c38c4c
44c6352c
63d0301c
0017311c
09c34664
0000931c
02930815
16c305c3
04bc29c3
0ef20b50
155c20e6
355c1e75
39840464
0467355c
d6bc05c3
00530b44
06961066
0f56e076
00000804
f9963016
217740c3
305c4137
40061e24
8000211c
6cd23283
0b44d6bc
60940007
1e24345c
0fdb303c
1e27345c
2d060b33
0b4d88bc
54940007
0444345c
0464245c
3f5cad00
3f5c00a1
2f5c00d5
2f5c0081
611700dd
13c7345c
245c4157
404713e7
345c0694
70721e24
1e27345c
202604c3
0b3eeabc
19540007
1e81245c
15544007
60376046
407742a6
60b76006
04c360f7
4d0615c3
01a03f3c
0b57debc
001c20c3
4007fec0
01f31d74
204605c3
34c342a6
0b4424bc
0050053c
01a01f3c
b0bc4046
40e608cb
0464345c
345c6d00
345c0467
7f721e24
1e27345c
d6bc04c3
07960b44
08040c56
40c33016
13c352c3
feb8201c
22946007
0b3eeabc
740c0cd2
1de4045c
201c6c00
20d7ff7c
30e401c3
740f15b4
1e24345c
0010341c
04c369f2
41462046
0b59c0bc
fec7201c
04c300f3
4c862026
0b59c0bc
02c320c3
08040c56
ff967016
42c360c3
606753c3
700c1435
700f6025
1fc30580
0b3f30bc
6065700c
6017700f
53e46085
06c30694
4e262046
0b59c0bc
feb8001c
0e560196
00000804
40c3f016
52c361c3
1dc4205c
305c340c
68f21e81
41462046
0b59c0bc
fe8b001c
305c0533
602715c9
305c0994
341c1e24
6bd22000
15a3005c
60470133
345c0694
010615c1
02946147
68200006
1de4045c
001c4c20
4007feb8
47d20d74
345c7880
245c0527
28800547
1de4745c
740f6780
0f560006
00000804
0336f016
40c3fc96
82c391c3
1404305c
feb9331c
72870354
40060494
1407245c
1e79345c
0c546147
c4bc04c3
00270ba3
345c0754
72871404
1fc67294
345c0e13
53c30464
1e546007
d6bc04c3
045c0b44
00071407
031c0a15
6194fecc
1e29345c
60076732
0b735b94
0604345c
05e4745c
58e4af80
301c07f4
345cff53
03c31407
58e409d3
28c34954
101c0aa0
bebc4000
145c0b3e
bebc47a3
60c30b3e
0660703c
17c304c3
0b4d88bc
2c940007
0444345c
0464245c
c0376d00
407742e6
00f700b7
13c304c3
79c327c3
debc7e80
00070b57
001c0415
0473fec0
0464345c
345c6c00
04c30467
0b44d6bc
0f150007
0607645c
05e7545c
fecc031c
345c0594
67321e29
045c6df2
01731407
345cb700
341c1e44
60070001
05c3b754
00060053
c0760496
08040f56
3f36f016
60c3f596
1e24305c
200603c3
6000111c
901c0183
00070000
0019c4dc
0003341c
07946047
01f7b0c3
02374066
04134277
0744065c
feb8901c
b2dc0007
60500018
00601b3c
3b3c2277
62370030
2dd21bc3
0784265c
484c4ad2
625741f7
62776d00
25002217
00732237
41f74006
365c40c6
df5c14c4
65d20124
65a02257
d2a4d3c3
47a3165c
22b725d2
4000131c
301c0435
62b74000
0000901c
31c32297
61b77f85
31c321d7
4d003b84
61374177
365c26f3
341c1e24
66d24000
801c79c3
c8c30005
365c03f3
6cf214c4
37c3e197
32e44157
72c30235
0090c73c
0009801c
0dc30153
bebc2297
70c30b3e
0050c03c
0005801c
202606c3
0b3eeabc
c21c03d2
06c30066
88bc1cc3
90c30b4d
34dc0007
365c0012
a3c30444
0464165c
365ca184
265c14c4
60071e24
32c35d94
4000341c
16946007
2f5c4166
c0770005
17c30ac3
625729c3
0b4464bc
202606c3
0b3eeabc
06c307f2
00501a3c
1abc4086
4ac30b51
02174884
f4bc14c3
06c30b3e
eabc2026
06f20b3e
14c306c3
1abc4066
821c0b51
d21c0003
ffa5fffd
20071bc3
4ac35354
0bc34884
f4bc14c3
06c30b3e
eabc2026
06f20b3e
14c306c3
1abc4066
06c30b51
eabc2026
00070b3e
000c84dc
0744365c
2c0c06c3
1abc2bc3
61d70b51
d2dc6007
365c000b
06c30784
41d72c0c
0b511abc
32c31693
4000341c
0ac367f2
42c617c3
24bc36c3
1bc30b44
1c542007
14c4565c
18345be4
0ea03bc3
bebc17c3
40c30b3e
0744365c
0ac36c0c
2e800884
b0bc24c3
848408cb
14c4365c
365c6e00
d4a414c7
41d7fe20
1d544007
1b54e007
14c4565c
0ea06117
bebc17c3
40c30b3e
0784365c
54a01bc3
0ac36c0c
2d000884
b0bc24c3
848408cb
14c4365c
365c6e00
d4a414c7
202606c3
0b3eeabc
44540007
ffb0583c
0415a007
ff7c901c
75c30cd3
1954a007
10f8101c
0000111c
8c0c640c
392c05c3
301c44c6
311c6590
46640017
04f270c3
ff83901c
1a3c0a13
25c30050
08cbb0bc
42c6a037
60264077
200660b7
06c320f7
2cc31ac3
debc37c3
c0c30b57
10f8201c
0000211c
8c4c680c
392c07c3
301c44c6
311c6590
46640017
0000c31c
9cc30315
365c0553
3c840464
0467365c
1e44365c
0008341c
06c365f2
0b44d6bc
1dc390c3
29c325d2
62dc4007
931cffec
1354feb9
165c2006
365c14c7
341c1e24
6bf20010
265c4066
00f31e6d
0003821c
fffdd21c
eab3ffa5
0b9609c3
0f56fc76
00000804
f096f016
305c40c3
341c1e24
a1861000
a48662f2
202604c3
0b8b08bc
000720c3
04c35a94
0096101c
0b4d88bc
000720c3
745c5294
645c0444
62860464
00053f5c
0f3c8077
15c30100
40bc35c3
345c0b44
341c1e24
66f20010
65a4201c
0017211c
201c00b3
211c65a0
04c30017
01401f3c
0b569ebc
000720c3
353c2e94
60370040
607762c6
60b76026
04c300f7
201c3f00
3f3c0096
debc0100
201c0b57
0007fec0
345c1a74
233c1e24
341c4004
43f20010
005369f2
614667d2
1e7d345c
345c6026
345c1e85
6c000464
0467345c
d6bc04c3
20c30b44
109602c3
08040f56
fb96f016
202640c3
0b3eeabc
ad8605d2
1e81245c
a0c642f2
15c304c3
0b4d88bc
000770c3
345c3b94
245c0444
cd000464
202606c3
34c34286
0b4424bc
78ad6026
202604c3
0b3eeabc
1a540007
1e81245c
16544007
01403f3c
233c4026
4026ffde
42864037
e0b74077
04c3e0f7
25c316c3
0b57debc
000750c3
70c30315
345c01f3
6e800464
0467345c
1e44345c
0008341c
04c365f2
0b44d6bc
07c370c3
0f560596
00000804
0f36f016
70c3f396
92c3b1c3
636463c3
0301005c
d2dc0007
875c000d
831c15c1
24540007
0007831c
831c09b4
0e540001
0004831c
000ce4dc
831c01f3
1c540008
0009831c
000c64dc
1eac0c53
9ebc36c3
80060aa1
301c1813
311c10fc
6c0c0000
1ecc8e8c
466436c3
1eec00b3
54bc36c3
40c30b1e
af3c1613
0ac301b0
41a62006
0891b0bc
202607c3
0b48dabc
01f01f3c
0b3f16bc
1501075c
011d0f5c
1509275c
01252f5c
1511375c
012d3f5c
075cbf06
742015b3
1f3c1980
08bc0260
4f3c0b3f
04c30280
3ac0173c
b0bc4086
0f3c08cb
19c302c0
b0bc28c3
275c08cb
3eec15b3
8037b520
60776186
09c37920
60b76180
af5c40f7
41a60087
01c34177
00801b3c
0080293c
fabc7700
09730b1d
01b08f3c
200608c3
b0bc41a6
07c30891
dabc2026
1f3c0b48
16bc01f0
275c0b3f
2f5c1501
375c011d
3f5c1509
075c0125
0f5c1511
bf06012d
15b3275c
19807520
02601f3c
0b3f08bc
02804f3c
173c04c3
40863ac0
08cbb0bc
02c00f3c
410619c3
08cbb0bc
15b3275c
b5203eec
61868037
79206077
618009c3
40f760b7
00878f5c
417741a6
1b3c01c3
293c0080
77000080
0a9d5ebc
800630c3
0f1534e4
1e24375c
4000341c
fecf401c
07c368f2
42862046
0b59c0bc
fecf401c
02800f3c
b8bc2186
00730b06
fec8401c
0d9604c3
0f56f076
00000804
0136f016
80c3e596
62c371c3
bcbc0fc3
a0060b1d
0fc300f3
26c317c3
0b1daabc
58e4a025
1b96f974
0f568076
00000804
0136f016
80c3cd96
62c371c3
5cbc0fc3
a0060b1d
0fc300f3
26c317c3
0b1d4abc
58e4a025
3396f974
0f568076
00000804
0136f016
80c3cd96
62c371c3
8cbc0fc3
a0060b1d
0fc300f3
26c317c3
0b1d7abc
58e4a025
3396f974
0f568076
00000804
00871016
00871954
002706d4
00470954
01932494
165400a7
1f9400c7
01c30333
23c312c3
0b5278bc
01c30313
23c312c3
0b537cbc
01c30253
23c312c3
0b5eacbc
01c30193
23c312c3
0b5ec4bc
01c300d3
23c312c3
0b5edcbc
08040856
005c26d2
680615d1
0b5ef4bc
00000804
0f36f016
70c3ec96
40b781c3
9f5c63c3
af5c03a4
6d0003c4
197439e4
00413f5c
201c13c3
2abc0100
4f3c0b49
96a40100
0007af5c
40774026
07c3be0c
28c314c3
566439c3
18c304c3
05d31984
00414f5c
409780f7
49c332e3
0680ae00
00613f5c
809713c3
402524c3
0b492abc
0100bf3c
1e540007
2f5c07c3
12c30061
00ff301c
4e208097
0b492abc
ab2029c3
0007af5c
60776026
07c39e0c
28c31bc3
466435c3
48c30bc3
26c33280
0b06c0bc
07c30573
00612f5c
301c12c3
809700ff
2abc4e20
b7200b49
0007af5c
40774026
07c39e0c
28c31bc3
466435c3
09c340c3
26c32097
0b493cbc
07c330c3
27c313c3
0b5f22bc
38c30bc3
26c32e80
0b06c0bc
04c303f2
001c83d2
1496fecf
0f56f076
00000804
0f36f016
70c3ed96
a3c391c3
15e9b05c
15c9305c
53946027
1e24405c
341c34c3
13c32000
105c63d2
08a015a3
640019c3
fff9335c
14c360b7
1000141c
00372dd2
0027af5c
19c307c3
3bc323c3
0b5f2abc
4f540007
3bc30c93
363cc9a0
81c3fff0
21c32097
053523e4
00478f5c
0001801c
3f5c07c3
13c30041
0100201c
0b492abc
78a02097
00c05f3c
fff0633c
0007af5c
40774026
07c39e0c
29c315c3
466436c3
05c340c3
2f0039c3
c0bc2bc3
00070b06
34c33494
600738a3
05f31c54
1b946007
c8a01bc3
00c05f3c
0007af5c
40774026
15c3820c
36c329c3
40c34664
39c305c3
2bc32f00
0b06c0bc
17940007
02b384d2
00732026
20b72006
15c9375c
06946047
15b3175c
2c0f6717
409700d3
3b846880
640f2717
00730006
fecf001c
f0761396
08040f56
3f36f016
50c3ff96
815c91c3
08c30003
4f540007
0014183c
4b942007
401cf42c
e007fe8d
d75c4854
41c30003
1cc306b3
29c36409
04892b00
03e40037
3bc32394
64a94c09
1e9423e4
14c305c3
0b4ae0bc
18540007
00011f5c
1e5d155c
3a84742c
255c4c89
05c31e65
0b8b34bc
000740c3
05c32294
1300193c
4c2b39c3
0b49a8bc
363c0353
63c30020
68e46364
343cd114
43c30020
4de44364
c0060c34
c33c7e00
a43c0040
2ac30010
b33c7d00
fdd30040
fe0b401c
019604c3
0f56fc76
00000804
0f36f016
40c3fb96
b2c371c3
0810a3c3
49dc6447
0f3c0013
28c30120
40462500
08cbb0bc
00993f5c
345c6077
00571569
13e410c3
001265dc
2b3403e4
1e24245c
2004323c
d2dc6007
345c0011
20571e89
30e401c3
001165dc
32c327f2
0b1b313c
0b5b313c
605700f3
002703c3
32c30a94
345c6d92
1f5c1e27
145c0021
0133156d
32c34057
05946047
00210f5c
156d045c
0020283c
033c704c
3d000300
b0bc4406
283c08cb
704c0220
135c3d22
104c0385
0381205c
05354407
105c2006
1bd30385
0230583c
13544007
0230323c
65dc3ae4
0a05000d
b0bc3e80
704c08cb
0381235c
345cb500
6b721e24
1e27345c
742008c3
3ae46065
000c35dc
0010353c
40b75da2
0010933c
345c7ea2
0f5c1e5d
045c0041
29c31e65
2fd23d22
1e24345c
011c0006
30830008
fe0a201c
02dc6007
131c000b
0d5400dd
1e24245c
000632c3
0008011c
65d23083
739232c3
1e27345c
0010593c
a40f1bc3
d52028c3
2e346ae4
eebc04c3
00070b95
363c2454
3ae40020
000875dc
1f3c1e80
3ebc00c0
593c0b3f
2f5c0030
18c30063
6e8068a0
78b43ae4
20372006
3e8004c3
68bc6006
20c30b95
76940007
00632f5c
0bc37500
0173600f
38843ac3
680f2bc3
345c00d3
6b921e44
1e47345c
345c6046
04c31e6d
eabc2006
07d20b3e
600c0bc3
1de4145c
600f6c80
48c4545c
1254a007
01403f3c
233c4606
04c3fc7e
11d0143c
345c23c3
566448e4
44940007
660760d7
345c4194
341c1e24
60070400
04c33054
0b4f90bc
25540007
34bc04c3
201c0b8b
0007fe0c
704c3194
2710033c
11d0143c
b0bc4606
345c08cb
341c1e24
1fe61000
04c364d2
0b9aa8bc
1e24345c
1000341c
04c364f2
0b858abc
145c20a6
01531e6d
1e24345c
0a9b303c
1e27345c
34bc04c3
20c30b8b
201c0133
00d3feb8
feba201c
201c0073
02c3fe78
f0760596
08040f56
50c3f016
02d261c3
701c24f2
34b3ff53
6025650c
002c600f
0084121c
0100201c
0892e6bc
4006742c
07fd235c
0ebc142c
03640892
0010303c
0867355c
1a84365c
21546007
1100053c
3500163c
b0bc4b86
301c08cb
311c10f8
6c0c0000
065c8c0c
155c1aa4
45462584
663c301c
0017311c
055c4664
07d20887
1a84165c
1aa4265c
08cbb0bc
0c67555c
0c84055c
1840163c
0100201c
0892e6bc
0c84355c
235c4006
055c07fd
0ebc0c84
03640892
0010303c
14c7355c
1d64365c
21546007
29c0053c
3ac0163c
b0bc4b86
301c08cb
311c10f8
6c0c0000
065c8c0c
155c1d84
45462584
663c301c
0017311c
055c4664
07d214e7
1d64165c
1d84265c
08cbb0bc
18c7555c
3200053c
2980163c
b0bc4406
365c08cb
355c15c4
5bcc18e7
00ff231c
053c0cd4
3bac3400
08cbb0bc
75005bcc
235c4006
00931a05
355c6006
065c1a05
240619e4
0b3ebebc
0ad220c3
2207055c
4440053c
19c4165c
08cbb0bc
055c0073
065c2207
24061a24
0b3ebebc
0ad220c3
2327055c
4680053c
1a04165c
08cbb0bc
055c0073
780c2327
20546007
0007182c
301c1d54
311c10f8
6c0c0000
155c8c0c
40c62584
663c301c
0017311c
055c4664
f06624c7
58ec0cd2
24a7255c
355c782c
380c24e7
b0bc582c
e00608cb
60077b8c
18ac2154
1e540007
10f8301c
0000311c
8c0c6c0c
2584155c
301c45a6
311c663c
46640017
2467055c
f06603f2
3b8c0173
b0bc58ac
58ac08cb
2487255c
355c78cc
053c2447
165c4a40
40061484
2584355c
0ba024bc
f06603d2
355c0153
0c0c2524
1444165c
1484265c
08cbb0bc
255c592c
60062547
1835365c
2544255c
2567255c
1819365c
25ad355c
1829265c
25c7255c
1843365c
25e6355c
1861265c
25f5255c
1869365c
25fd355c
1821265c
2605255c
1871365c
260d355c
1879265c
2615255c
1809365c
261d355c
1881265c
2625255c
1924365c
22546007
1944065c
1e540007
10f8301c
0000311c
8c0c6c0c
2584155c
301c4666
311c663c
46640017
2647055c
f06603f2
165c0173
265c1924
b0bc1944
365c08cb
355c1944
265c2667
255c1761
365c2685
355c1891
365c268d
60071964
065c2254
00071984
301c1e54
311c10f8
6c0c0000
155c8c0c
46662584
663c301c
0017311c
055c4664
03f226a7
0173f066
1964165c
1984265c
08cbb0bc
1984265c
26c7255c
1839365c
26e5355c
1899265c
26ed255c
19a4365c
2507355c
0f5607c3
00000804
3f36f016
50c3e896
c2c391c3
081043c3
49dc6047
01c3002d
1f3c0884
30bc05c0
2cc30b3f
6065680c
45d7680f
ff7c601c
4000231c
002ce5dc
ed0038a4
e4dc74e4
4f3c002b
40060140
af3c40f7
06930580
03c360d7
04940127
fe90601c
1cc35753
323c440c
38a40030
85dc37e4
19c3002a
1ac30500
0b3f30bc
680c2cc3
0030233c
4c0f3cc3
08c32597
6c806820
65dc37e4
300f0029
610009c3
ffe7345c
1cc36880
65d7640f
45977fa5
65f76d20
03c360d7
00f70025
c5d78105
cb94c007
10f8301c
0000311c
8c0c6c0c
0408001c
44c616c3
6604301c
0017311c
70c34664
12dc0007
203c0027
40772d80
631260d7
06000f3c
b33c6180
af5cfac0
c0370064
a21c11d3
1bc3ffff
d15c2410
07c3ffe4
29c31dc3
fcbc752c
355c0ab0
361c1e24
940c0040
200607c3
098b233c
56bc718c
40c30ac2
1e24355c
0404833c
400728c3
7cec1d94
0206331c
331c0f54
16940285
1ed2255c
c3dc4007
23640023
32e47c2c
002370dc
255c0173
40071ee2
0022e3dc
7c2c2364
90dc32e4
80070022
175c4694
20071819
28c33354
30944007
0d8c740c
34bc2057
00070ba7
8f5c2994
0f3c02c7
19c30580
752c4086
0ba024bc
000760c3
301c0a15
311c10f8
6c0c0000
07c38c4c
3ef318c3
0c0c6597
29c31dc3
08cbb0bc
0d8c740c
05801f3c
34c34046
0ba83abc
c02760c3
c0070354
740c1194
135c6d8c
2bd202b1
02b9235c
0dac48d2
400617c3
0b9f7abc
005360c3
c4d264c3
62f26017
07c3c037
0aa364bc
fff8b21c
0001a31c
fff716dc
1ac39ac3
32dc2007
07c30013
41572117
fcbc752c
355c0ab0
361c1e24
940c0040
200607c3
098b233c
56bc718c
60c30ac2
031c06d2
0f54ff74
6dd2750c
6d8c740c
02b1035c
0dac0bd2
400617c3
0b9f7abc
009360c3
20b72026
40060073
053c40b7
17c34080
0b61eebc
706730c3
20970454
15542007
64bc07c3
301c0aa3
311c10f8
6c0c0000
07c38c4c
44c62006
6604301c
0017311c
655c4664
31731407
1e24355c
355c7b72
801c1e27
811c10f8
28c30000
8c0c680c
0100001c
44c62097
6604301c
0017311c
90c34664
07c30af2
0aa364bc
600c08c3
07c38c4c
1d532097
231c5fcc
0ad400ff
b0bc3fac
7fcc08cb
00410f5c
09a129c3
2f5c00b3
19c30041
355c440d
341c1e24
60070040
255c1194
4ed204e4
3fcc1fac
0b472ebc
07c309f2
04e4155c
0b5590bc
601c03f2
7cecfebe
0206331c
331c5054
84dc0285
40060009
055c45b7
00071f44
301c1494
311c10f8
6c0c0000
001c8c0c
352c0098
301c4146
311c6604
46640017
1f47055c
0f930cf2
1f61355c
e6bc6fd2
00060b1c
1f65055c
1f44055c
255c352c
e6bc4764
00070b0e
1c0c6b94
05801f3c
1f44255c
42bc7c2c
00070ac0
20266194
1f65155c
5e94c007
1e24355c
0040341c
58946007
1f44055c
0b1c4cbc
355c20c3
23e41ed2
601c4f15
0993fe67
1fa4055c
13940007
10f8301c
0000311c
8c0c6c0c
352c0a06
301c44a6
311c6604
46640017
1fa7055c
1a730cf2
2019155c
b6bc2dd2
40060ad2
201d255c
1fa4055c
255c352c
5ebc4764
1cec0ace
21c32006
0ace82bc
1c0c30c3
255c3c2c
d6bc1fa4
00070acf
60261794
201d355c
1494c007
1e24355c
0040341c
055c6ff2
72bc1fa4
20c30ace
1ee2355c
061523e4
fe66601c
601c0073
07c3feaa
0aa364bc
10f8801c
0000811c
640c18c3
07c38c4c
44c62006
6604301c
0017311c
28c34664
8c0c680c
20060406
301c44c6
311c6604
46640017
0df270c3
600c08c3
09c38c4c
44c617c3
6604301c
0017311c
0e734664
24d22017
61c3c3f2
c0070073
355c2d54
341c1e24
60070040
363c2594
85460970
02b46027
750c85a6
12546007
60d7dcaf
00067ccf
3c511cef
3c8f34ec
4080353c
750c7c2f
366417c3
c00603d2
05c30173
24c32046
0b59c0bc
1e24355c
355c7072
655c1e27
355c1407
341c1e24
69d20040
16a0363c
05b46027
355c6006
00531407
355ccbf2
341c1e24
63c30010
006665d2
1e6d055c
05c3c006
eabc2006
07d20b3e
640c1cc3
1de4255c
640f6d00
10f8501c
0000511c
8c4c740c
200607c3
301c44c6
311c6604
46640017
8c4c740c
200609c3
301c44c6
311c6604
46640017
601c0193
0133feb8
00f3d066
fe66601c
601cc3f3
c393fe67
189606c3
0f56fc76
00000804
1f36f016
40c39e96
b2c391c3
e80c83c3
b9dc6447
0f3c001d
27801860
b0bc4046
1f5c08cb
145c0c33
145c1576
31c31e24
4000341c
1569245c
3f5c66f2
23e40c39
0d5310b4
00ff231c
231c6754
645400fd
0c393f5c
00ff331c
331c5f54
5c5400fd
2004313c
42dc6007
1f5c001b
22770c39
1e89345c
c5dc31e4
6257001a
345c6ff2
02571e24
0b1b303c
0b5b303c
1e27345c
01212f5c
156d245c
62570313
c31cc3c3
0b940001
1e24345c
345c6d92
0f5c1e27
045c0121
0133156d
21c32257
05944047
01213f5c
156d345c
1563045c
01660f5c
345c302c
233c1e24
2f5c0d8b
233c0006
2f5c0dcb
233c0026
2f5c0e4b
233c0046
2f5c0d4b
233c0066
2f5c0e8b
333c0086
3264090b
01c36177
02c01f3c
60064026
0b400ebc
245c0113
3f5c1569
23e40c39
001570dc
0020273c
033c704c
39c30100
44062d00
08cbb0bc
0220373c
61a209c3
573c6237
a01c0230
7fe50000
3f5c61f7
63c700e1
a01c03b4
62170001
c31cc3c3
04540020
00070ac3
22171c54
646531c3
b5dc38e4
704c0012
0500033c
2e8039c3
b0bc4217
704c08cb
01010f5c
0385035c
b4802217
1e24345c
345c6a72
00b31e27
40074217
001124dc
604577a0
d5dc38e4
19c30010
1f3c0680
3ebc0300
a0450b3f
01832f5c
0010323c
6e806fa0
d5dc38e4
231c000f
95dc012c
0f3c000f
39c30340
b0bc2e80
0f5c08cb
74000183
1f5c2006
09c30196
28094180
033c22b7
51c30010
6c8063a0
15dc38e4
2007000e
000e42dc
61c32006
63f26829
00b32026
00dd331c
c0260294
c3c36297
ffffc21c
00c7cf5c
00c13f5c
402562b7
ed946007
345cb400
00061e24
0008011c
0f5c3083
20c30141
402622d2
63f22264
10944007
7f3233c4
ccf262d2
72dc6007
4007000b
000b42dc
1e24345c
345c7392
1bc31e27
d7a0a40f
363468e4
eebc04c3
00070b95
04c32d54
f8bc2026
00070b93
000a04dc
0020363c
35dc38e4
19c30009
1f3c0680
3ebc1840
a0450b3f
0c232f5c
6e806ba0
55dc38e4
3f3c0008
60370300
39c304c3
60262e80
0b9568bc
14dc0007
0f5c0008
74000c23
640f1bc3
28c300b3
0bc36b80
20e6600f
1e75145c
1e24345c
345c6b72
341c1e27
60070400
704c5c54
133c04c3
40262710
0ba07cbc
1e44245c
2004323c
043c64d2
00f30f40
65d23ac3
4004323c
4d546007
005c0fd2
345c02d3
63321e49
0001341c
125430e4
8004323c
60070af2
345c3854
303c1e24
345c0a9b
06331e27
fe62001c
2d946007
04c30753
03001f3c
0b6044bc
001c30c3
6007fe0c
704c3074
133c10cc
44060300
0b1bf6bc
400720c3
345c2694
341c1e24
65d21000
a8bc04c3
20c30b9a
1e24345c
1000341c
04c365f2
0b858abc
610620c3
1e75345c
01f302c3
1f3c04c3
44bc0300
01330b60
feb8001c
001c00d3
0073feba
fe0a001c
f8766296
08040f56
60c37016
03e1305c
200664d2
0b4e4abc
10f8501c
0000511c
8c4c740c
392c182c
301c43c6
311c66a4
46640017
782f6006
8c4c740c
392c186c
301c45c6
311c66a4
46640017
786f6006
15c9365c
365c67d2
341c1e24
60072000
365c1f94
341c1e44
60070040
18cc1954
0b1c08bc
10f8301c
0000311c
8c4c6c0c
392c18cc
301c4406
311c66a4
46640017
78cf6006
1e44365c
365c6692
365c1e47
341c1e44
65d20020
202606c3
0b54ecbc
1f44065c
15540007
0b1ce6bc
10f8301c
0000311c
8c4c6c0c
1f44065c
4146392c
66a4301c
0017311c
60064664
1f47365c
1f84065c
1b540007
2011365c
b6bc66d2
60060ad2
2015365c
10f8301c
0000311c
8c4c6c0c
1f84065c
44a6392c
66a4301c
0017311c
60064664
1f87365c
1fa4065c
1b540007
2019365c
b6bc66d2
60060ad2
201d365c
10f8301c
0000311c
8c4c6c0c
1fa4065c
44a6392c
66a4301c
0017311c
60064664
1fa7365c
1fc4065c
1b540007
2021365c
b6bc66d2
60060ad2
2025365c
10f8301c
0000311c
8c4c6c0c
1fc4065c
44a6392c
66a4301c
0017311c
60064664
1fc7365c
0704065c
165c05d2
b8bc0724
501c0b06
511c10f8
740c0000
065c8c4c
392c0704
301c41e6
311c66a4
46640017
365c6006
740c0707
065c8c4c
392c06c4
301c41e6
311c66a4
46640017
365c6006
365c06c7
67f20639
1e24365c
0010341c
21546007
10f8501c
0000511c
8c4c740c
0684065c
41e6392c
66a4301c
0017311c
60064664
0687365c
8c4c740c
0644065c
41e6392c
66a4301c
0017311c
60064664
0647365c
0abc06c3
365c0ba8
60071371
301c1a54
311c10f8
6c0c0000
065c8c4c
392c0b44
301c4726
311c66a4
46640017
16e0363c
0b47365c
365c6006
60061375
0b66365c
08040e56
3f36f016
40c3bd96
d2c32037
b3d7a3c3
15e9805c
15f1b05c
14bc15c3
90c30ba0
1010cf3c
20060cc3
b0bc4106
6f3c0891
2f5c10c0
263c09c1
0ac3fede
10a01f3c
0b3f08bc
15c304c3
0b48dabc
10501f3c
0b3f16bc
15d1345c
40946027
06404f3c
eebc04c3
04c30b00
28c319c3
0b05a6bc
101c04c3
111c6330
2bc30017
0b05a6bc
1cc304c3
a6bc4106
04c30b05
406616c3
0b05a6bc
1dc304c3
a6bc2ac3
5f3c0b05
04c30c10
5cbc15c3
04c30b05
28c319c3
0b05a6bc
101c04c3
111c6360
2bc30017
0b05a6bc
15c304c3
a6bc28c3
04c30b05
5cbc2017
e0060b05
5f3c0833
05c30040
0b1decbc
000770c3
05c33994
28c319c3
0b1ddabc
101c05c3
111c6330
2bc30017
0b1ddabc
1cc305c3
dabc4106
05c30b1d
406616c3
0b1ddabc
1dc305c3
dabc2ac3
4f3c0b1d
05c30c10
cabc14c3
05c30b1d
28c319c3
0b1ddabc
101c05c3
111c6360
2bc30017
0b1ddabc
14c305c3
dabc28c3
05c30b1d
cabc2017
07c30b1d
fc764396
08040f56
f896f016
41c350c3
b2dc0007
20070013
001382dc
6007602c
001342dc
715c000c
03d20361
0bae02bc
0080643c
cabc06c3
72c60b23
c4dc0007
706c0012
706f6025
ccbc06c3
940f0b23
4c0b700c
1566255c
0323345c
2006355c
255c534c
730c1fe7
14a7355c
550f52ec
355c500c
48491e24
091b323c
1e27355c
13c3500c
133c6869
155c0a5b
345c1e27
355c0261
313c1e8d
68f20104
245c31c3
323c0229
355c0d9b
355c1e27
245c1e24
323c0231
355c0ddb
245c1e27
323c0239
355c0e5b
245c1e27
323c0221
355c0d5b
23c31e27
0241345c
0e9b233c
1e27255c
1e44055c
0361345c
09db033c
1e47055c
0273345c
1eb6355c
0283345c
1ed6355c
0293345c
1ee6355c
245c32c3
323c0201
355c089b
245c1e27
323c0209
355c08db
245c1e27
323c01e1
355c095b
245c1e27
323c01e9
355c099b
245c1e27
323c01f1
355c09db
245c1e27
323c01f9
355c0a1b
13c31e27
0211345c
101b133c
1e27155c
245c30c3
323c0249
355c081b
245c1e47
323c0251
355c085b
245c1e47
323c0259
355c08db
313c1e47
6df20104
255c50ac
70cc0647
0667355c
255c50ec
710c0687
06a7355c
255c512c
714c0747
0787355c
255c516c
91ac0767
142c81b7
14c387d2
0154201c
08cbe6bc
3f5c0113
13c300c1
0154201c
0891b0bc
1e24255c
0104423c
355c142c
1f3c1563
800701c0
3f5c1e94
323c00e6
3f5c0d8b
323c0006
3f5c0dcb
323c0026
3f5c0e4b
323c0046
3f5c0d4b
323c0066
3f5c0e8b
323c0086
3264090b
40266177
039334c3
00e63f5c
3f5c6026
323c0006
3f5c0dcb
323c0026
3f5c0e4b
323c0046
3f5c0d4b
323c0066
3f5c0e8b
323c0086
3264090b
40266177
0ebc6006
355c0b40
341c1e24
60070010
e0071494
355c1294
6cd20744
6ad26c0c
0764055c
600c07d2
009368f2
ff53301c
301c00b3
0053fec3
03c36026
0f560896
00000804
ff96f016
71c350c3
201c2006
b0bc0920
5dcc0891
353c552f
776f0640
37cf20a6
0800353c
0447355c
04a7155c
4080053c
a0bc2006
5fe60b4e
1427255c
1447255c
355c6006
355c4827
355c48a7
355c4887
355c4847
101c4867
74800904
74af748f
255c4006
255c1e6d
255c1e75
255c1e95
255c1e9d
255c1e7d
301c1e55
311cd368
760f0016
101cb5ef
155c4000
5fe647a6
1387255c
13a7255c
13c7255c
13e7255c
68bc05c3
053c0b3f
aabc2b00
601c0b3f
611c10f8
780c0000
001c8c0c
352c02a4
301c4426
311c66dc
46640017
0007144f
000872dc
201c2006
b0bc02a4
780c0891
001c8c0c
352c0154
301c43c6
311c66dc
46640017
0007142f
05c37354
66bc17c3
00370b6a
202710c3
40066d94
1561355c
00fe331c
3f5c0494
23c30001
1e24355c
0b9b323c
1e27355c
10f8601c
0000611c
8c0c780c
0428001c
45c6352c
66dc301c
0017311c
146f4664
4a540007
01c8021c
0b00eebc
033c746c
ecbc1680
00370b1d
40940007
033c746c
bcbc2240
00370b1d
38940007
033c746c
5cbc2900
00370b1d
30940007
033c746c
8cbc35c0
00370b1d
28940007
74cf7c2c
17946007
8c0c780c
352c0206
301c4406
311c66dc
46640017
000714cf
355c1554
66721e44
1e47355c
0b1c16bc
0ef20037
155c2006
155c48c7
353c48e7
355c16e0
20370b47
50660073
00174037
0f560196
00000804
0736f016
80c3f496
52c341c3
af5c60f7
9f5c02a4
c5d702c4
01007f3c
98bc07c3
45170aca
07c34037
25c314c3
d4bc60d7
40c30aca
cdd20ef2
68cc28c3
4617c037
07c34077
2ac313c3
0cbc39c3
40c30acc
10948007
6c0c39c3
46576037
66974077
0f3c60b7
26d70100
3ac34717
0acb28bc
0f3c40c3
1ebc0100
04c30acb
e0760c96
08040f56
0136f016
80c3f696
52c341c3
7f3c63c3
07c30080
0aca98bc
40374417
14c307c3
36c325c3
0acad4bc
0ef240c3
68cc28c3
403744d7
40774517
13c307c3
64974457
0acc0cbc
0f3c40c3
1ebc0080
04c30acb
80760a96
08040f56
41c31016
105c44f2
00732003
2c0c684c
24c300cc
0adcb2bc
08040856
12c301c3
605723c3
0adcb6bc
00000804
0f3cfd96
00370080
00770157
12c301c3
611723c3
0adef4bc
609703f2
001c63f2
0396feb6
00000804
fe961016
803780cc
00770157
12c301c3
611723c3
0adc6abc
08560296
00000804
fe967016
940ca197
c037c1d7
c077c0cc
12c301c3
34c323c3
0b1cccbc
03f40007
0006140f
0e560296
00000804
1f36f016
60c3f596
42b74006
60064277
1ea5305c
15d9305c
12546047
20546107
fe8a501c
0000b01c
04dc6027
305c001f
60071f44
001e12dc
1f61305c
305c01b3
60070644
001d92dc
0684305c
42dc6007
305c001d
a00606c4
46946007
205c39b3
4cd215f9
1fa4705c
62dce007
305c001c
60072019
001c12dc
705c0173
e0071f84
001bb2dc
2011205c
62dc4007
7c4c001b
22dc6007
301c001b
311c10f8
6c0c0000
0a068c0c
44a6392c
63b8301c
0017311c
198f4664
b0c3b066
82dc0007
64a6001a
392c79af
4764265c
0ace5ebc
000750c3
001994dc
398c06c3
16bc27c3
50c30b6d
04dc0007
40260019
1ea5265c
0200301c
701c6277
711c10f8
7c0c0000
001c8c0c
20060200
301c44c6
311c63b8
46640017
0007b0c3
0017a2dc
15d9365c
1f546047
31546107
b4dc6027
784c0016
133c18cc
46060710
0b1bf6bc
000750c3
001674dc
265c784c
235c1571
784c038d
1579265c
0395235c
4606784c
06934c2f
0200301c
0587365c
8c0c7c0c
0200001c
44c62006
63b8301c
0017311c
065c4664
00070567
28731e94
02c03f3c
0200201c
fe7e233c
1b3c198c
23c30010
0ad14cbc
fe9e501c
44dc0007
2f5c0013
3bc30141
62974c0d
62776025
0200301c
009362b7
64dca007
40460012
1ea5265c
15d9365c
19546047
3e546107
34dc6027
584c0011
02403f3c
365c6037
60771f44
60b76006
613760f7
123c06c3
46060710
50bc3bc3
07930b6d
165c584c
465c0644
565c0664
365c0684
603706a4
0564365c
363c6077
60b70b00
0067bf5c
02403f3c
365c6137
617706c4
06e4365c
323c61b7
61f70710
0040323c
06c36237
35c324c3
0b6ca8bc
265c02b3
44d215f9
1fa4565c
565c0073
798c1f84
2f3c984c
40370280
13c306c3
343c25c3
24bc0710
50c30b6d
84dc0007
6066000c
1ea5365c
15d9365c
92dc6007
6047000b
61070735
000b44dc
4297784c
60864c2f
1ea5365c
1e24165c
1000141c
365c26f2
71c315d9
02946047
365ce046
610715d9
60a70554
60c70354
e0060294
7d004257
0090933c
202606c3
0b3eeabc
921c03d2
06c30066
88bc19c3
50c30b4d
e4dc0007
365c0008
a3c30444
0464265c
0ac3a284
3d806257
36c34206
0b444abc
e8d28126
01230f5c
00901a3c
0b3f08bc
2ac38166
1bc30a00
b0bc4257
e25708cb
202606c3
0b3eeabc
000730c3
373c3954
ee00ffb0
10f8c01c
0000c11c
680c2cc3
07c38c0c
44c6392c
63b8301c
0017311c
80c34664
53540007
00501a3c
b0bc27c3
e03708cb
607762c6
40b74026
60f76006
1ac306c3
38c329c3
0b57debc
2cc390c3
8c4c680c
392c08c3
301c44c6
311c63b8
46640017
0000931c
59c30b15
06c30633
29c31ac3
0b5004bc
000750c3
40a62994
1ea5265c
0464365c
365c3984
365c0467
341c1e44
65f20008
d6bc06c3
50c30b44
531ca4d2
1494feb9
4ebc06c3
02d20b88
410650c3
1e75265c
501c0173
0093fec4
fe8a501c
b01c00b3
00530000
784cb066
0710033c
b8bc2c2c
784c0b06
4c2f4006
6fd23bc3
10f8301c
0000311c
8c4c6c0c
392c0bc3
301c44c6
311c63b8
46640017
7ebc06c3
05c30b51
f8760b96
08040f56
12c301c3
609723c3
0b1cb8bc
04f40007
0c0f6057
08040006
1f36f016
60c3f496
c2c3b1c3
2810a3c3
22b72006
205c4006
205c1ea5
323c1e24
9fe60104
f4dc6007
305c001f
60c71e71
204608b4
c0bc4146
401c0b59
3e73fe8b
0a04323c
00a0331c
32c30b94
111c2006
31830800
fea7401c
52dc6007
323c001e
331c1204
0b940120
200632c3
2800111c
401c3183
6007fea7
001e22dc
15d9365c
16546047
0a546107
34dc6027
365c001c
6c0c0764
fec3401c
265c0113
48f215f9
fe9f401c
2021365c
d2dc6007
0026001b
1ea5065c
15d9365c
72dc6047
6107000f
60276554
001a64dc
22772006
10f8301c
0000311c
8c0c6c0c
0098001c
4146392c
6614301c
0017311c
198f4664
42dc0007
41460019
392c59af
4764265c
0b0ee6bc
000740c3
001904dc
0764365c
1f3c0c0c
598c0240
b4bc6c4c
40c30abe
34dc0007
198c0018
0b1c4cbc
40c350c3
b3dc0007
365c0017
401c1ed2
53e4fe67
001743dc
784c85c3
2c2f2606
1e24365c
1000341c
600779c3
a31c1254
09dc0001
0bc30016
1f3c0984
3ebc02e0
3f5c0b3f
35e40173
001584dc
0020793c
74a019c3
3ae46f80
0014d5dc
62b76006
765c14d3
365c1fc4
43c315f9
37546007
02770006
10f8301c
0000311c
8c0c6c0c
392c0a06
301c44a6
311c6614
46640017
0007198f
0012d2dc
39af24a6
265c392c
5ebc4764
40c30ace
94dc0007
365c0012
0c0c0764
02401f3c
6c4c598c
0ab1a4bc
0df240c3
07c3f98c
0ace72bc
365c20c3
23e41ee2
401c0415
2233fe66
20071ac3
001092dc
39c32bc3
309d823c
0010383c
05dc3ae4
065c0010
00071f84
301c1394
311c10f8
6c0c0000
0a068c0c
44a6392c
6614301c
0017311c
065c4664
0df21f87
165c1cf3
20072011
b6bc1154
40060ad2
2015265c
1f84065c
265c392c
5ebc4764
40c30ace
b4dc0007
593c000d
7c4c0010
06801bc3
265c18c3
6c2c1f84
0acfd6bc
401c04d2
1973fea0
265c4026
301c2015
79cf0200
34dc8007
08c3000c
02f3e280
0001a31c
000b79dc
09840bc3
02e01f3c
0b3f3ebc
01732f5c
0020323c
a5dc3ae4
793c000a
59cf0020
0000801c
165c2046
365c1ea5
604715d9
61072b54
60271654
000944dc
0380363c
598c6037
60064077
60f760b7
06c36137
2b802bc3
3f3c28c3
8cbc0280
06f30b6f
1fc4165c
15f9365c
398c62d2
1f84365c
263c984c
40370380
23c306c3
0710343c
0b6d24bc
584c0493
0644165c
0664465c
0684565c
06a4065c
365c0037
60770704
0e40363c
000660b7
013700f7
63800bc3
7b8b6177
323c61b7
61f70710
0040323c
06c36237
35c324c3
0b6ca8bc
000740c3
00665294
1ea5065c
15d9365c
20546047
1a546107
3d946027
460759cc
22974294
3f542007
033c784c
b0bc0710
784c08cb
233c6f8c
365c820b
401c1573
23e4febb
78843294
784c00f3
2c2f39cc
5b8b0073
6086fd00
1ea5365c
4ebc06c3
40c30b88
21940007
065c00a6
1cc31ea5
4106e40f
1e75265c
1e24365c
0020341c
13546007
06c3786c
0b40133c
0b5408bc
017340c3
fe8a401c
90660113
401c00d3
0073feb8
fec2401c
033c784c
2c2c0710
0b06b8bc
0006784c
06c30c2f
0b517ebc
0c9604c3
0f56f876
00000804
ff963016
12c301c3
a15743c3
22540007
20546007
1e54a007
ff7c201c
0200131c
3f3c1eb4
40060040
fe7e233c
35c32fc3
0b1c72bc
000720c3
211712f4
03e431c3
20170c94
04c32ad2
08cbeabc
07d220c3
201c0093
0073ff53
fe6d201c
019602c3
08040c56
12c301c3
605723c3
0b1c72bc
00000804
3f36f016
60c3f796
417791c3
0006b3c3
01160f5c
20064810
d65c21f7
400615e1
1ea5265c
15d9765c
0754e047
fe8a501c
64dce107
13f30030
0001b31c
002fc9dc
02208f3c
0a8409c3
3ebc18c3
0f5c0b3f
303c0113
3be40020
002ee5dc
1eb3365c
093530e4
17c306c3
c0bc4506
501c0b59
5cd3fe6f
10f8c01c
0000c11c
640c1cc3
392c8c0c
301c41e6
311c65e0
46640017
0647065c
22dc0007
4a3c002d
2f5c0020
265c0113
39c30667
b0bc2e00
3f5c08cb
91800113
1ec6365c
7e007aa4
b5dc3be4
19c3002b
18c30600
0b3f3ebc
0020543c
01130f5c
61202ac3
3be46e80
002ac5dc
680c2cc3
392c8c0c
301c41e6
311c65e0
46640017
0687065c
02dc0007
3f5c002a
365c0113
29c306a7
23c32a80
08cbb0bc
01133f5c
7e009580
d5dc3be4
19c30028
18c30600
0b3f3ebc
0020543c
01130f5c
61202ac3
3be46e80
0027e5dc
6c0c3cc3
392c8c0c
301c41e6
311c65e0
46640017
06c7065c
22dc0007
2f5c0027
265c0113
39c306e7
b0bc2e80
85c308cb
01130f5c
0d938084
0003b31c
0025e9dc
0ac329c3
501c6822
6067fea2
0025b4dc
00203a3c
09a229c3
0b4a90bc
501c80c3
0007fea1
0024f3dc
00307a3c
63a209c3
01163f5c
3be46085
002405dc
1f84065c
13940007
10f8301c
0000311c
8c0c6c0c
392c0a06
301c44a6
311c65e0
46640017
1f87065c
44f30ef2
2011365c
600753c3
b6bc1154
40060ad2
2015265c
1f84065c
265c392c
5ebc4764
50c30ace
a4dc0007
473c0021
08c30010
21c32006
0ace82bc
19c330c3
1f5c0600
265c0113
d6bc1f84
04d20acf
fea0501c
3f5c40b3
40260113
2015265c
e4dca007
84c3001f
20268384
1ea5165c
15d9365c
07b460c7
51dc6087
6047000d
00d30494
04546107
fe8a501c
365c3d33
00061e24
4000011c
60073083
000c44dc
3aa438c3
c364c3c3
040cc31c
001d45dc
d2bc06c3
00070b3e
08c32354
3aa438c3
3be46045
001c85dc
0010283c
d33c39c3
6c22209d
10546087
04b46087
09946047
60a701b3
60c70454
35930494
3573a0c6
ff7b501c
a0a61553
a08634d3
a1063493
0001d31c
a0860254
cebc05c3
01b70b23
3aa438c3
3be46045
0019e5dc
088409c3
02201f3c
0b3f3ebc
0002821c
01132f5c
3aa432c3
3be43884
0018e5dc
04007c3c
10f8b01c
0000b11c
640c1bc3
07c38c0c
44c6392c
65e0301c
0017311c
065c4664
00070567
001762dc
0587765c
f0bc05c3
065c0b23
2bc305c7
8c0c680c
44c6392c
65e0301c
0017311c
065c4664
000705a7
001602dc
065c784c
133c0564
44060100
08cbb0bc
0564365c
033c584c
123c0200
44060300
08cbb0bc
0564365c
0400033c
1a8419c3
b0bc2cc3
365c08cb
265c0564
465c0584
065c05a4
003705c4
13c305c3
7cbc34c3
50c30b25
a4dc0007
d31c0013
08540001
ff7b501c
0003d31c
001314dc
365c0193
60071f44
001212dc
1f61365c
c2dc6007
01330011
2019065c
62dc0007
00730011
21b72006
265c4046
365c1ea5
60c715d9
608706b4
60476634
01130494
06546107
fe8a501c
0000a01c
765c1d33
20061e24
4000111c
e0077183
301c5494
311c10f8
6c0c0000
0f5c8c0c
392c0113
301c44c6
311c65e0
46640017
0007a0c3
000e82dc
188419c3
01132f5c
08cbb0bc
0001d31c
501c0854
d31cff7b
04dc0003
0313000c
01133f5c
1f44165c
e0772037
e0f7e0b7
1ac306c3
3f3c23c3
eebc01c0
50c30b71
f3dc0007
90c3000a
57c39364
3f5c03b3
465c0113
065c05a4
003705c4
1fa4165c
e0b72077
e137e0f7
1ac306c3
34c323c3
0b6d2cbc
90c350c3
34dc0007
00930009
95c3a006
4066a5c3
1ea5265c
15d9365c
06b460c7
6b346087
04946047
610700d3
501c0454
0f53fe8a
1e24365c
111c2006
31834000
5b946007
01132f5c
d31c8284
07540001
ff7b501c
0003d31c
09f36794
d2bc06c3
00070b3e
301c3d54
311c10f8
6c0c0000
001c8c0c
392c0200
301c44c6
311c65e0
46640017
03f270c3
09d3b066
05a4165c
05c4265c
94bc6197
09e40ab5
81d70e94
101c8cd2
bebc0200
30c30b3e
17c304c3
eabc23c3
03d208cb
feb6501c
10f8301c
0000311c
8c4c6c0c
392c07c3
301c44c6
311c65e0
46640017
2694a007
931c01d3
20940024
000701d7
165c1d54
29c305a4
08cbeabc
16940007
365c6086
06c31ea5
eabc2006
04d20b3e
1de4065c
20a68084
1ea5165c
08114157
365c6086
a0061e6d
501c0073
0ac3feb6
1e540007
10f8301c
0000311c
8c4c6c0c
392c0ac3
301c44c6
311c65e0
46640017
a0e601f3
0010823c
501ccc13
0113fec4
00d3b066
feb8501c
501c0073
06c3fed1
0b517ebc
099605c3
0f56fc76
00000804
1f36f016
50c3f996
c2c3a1c3
200673c3
40062177
00d62f5c
cc0c3cc3
105c2026
d2bc1ea5
46c30b3e
0002801c
e02709d2
0012c9dc
833c3ac3
463c609d
73200020
37e46045
001225dc
0a002ac3
01a01f3c
0b3f3ebc
0020b43c
00d32f5c
3b846b20
35dc37e4
231c0011
f5dc0200
155c0010
20072019
946c2e54
0c40343c
05a7355c
255c4286
05c305c7
0b3ed2bc
21540007
0004831c
343c0994
355c0d80
240605a7
05c7155c
831c02d3
09940005
0f80343c
05a7355c
355c6606
017305c7
0006831c
343c0894
355c1280
480605a7
05c7255c
355c6046
255c1ea5
40071f44
155c1c54
20071f61
3f5c1854
403700d3
40774006
40f740b7
1ac305c3
23c31b84
01403f3c
0b71eebc
901c60c3
09e40000
90c30674
0073c006
96c3c006
2019155c
17542007
00d33f5c
05a4455c
05c4255c
155c4037
20771fa4
40b74006
413740f7
1ac305c3
23c31b84
2cbc34c3
60c30b6d
f4dcc007
60660009
1ea5355c
1f44355c
62dc6007
155c0008
20071f61
000812dc
d2bc05c3
00070b3e
746c6d54
00c4321c
05a7355c
255c4286
301c05c7
311c10f8
6c0c0000
001c8c0c
16c30200
301c44c6
311c6628
46640017
03f270c3
0e33d066
0005831c
831c1354
1b540006
831c6b06
21940004
321c746c
355c00d8
640605a7
05c7355c
019e301c
746c02d3
00f8321c
05a7355c
155c2606
301c05c7
0173019f
321c746c
355c0128
480605a7
05c7255c
01a0301c
155c07c3
255c05a4
94bc05c4
90e40ab5
81570e94
101c8cd2
bebc0200
30c30b3e
17c304c3
eabc23c3
03d208cb
feb7601c
10f8301c
0000311c
8c4c6c0c
200607c3
301c44c6
311c6628
46640017
931c01f3
0a940024
08d20157
133c746c
29c30b40
08cbeabc
601c03d2
355cfeb7
7c721e24
1e27355c
2f5c1bc3
650000d3
640f1cc3
255c40a6
00731ea5
feb8601c
355c6006
355c05a7
05c305c7
0b517ebc
079606c3
0f56f876
00000804
0336f016
40c3fc96
52c361c3
8f5ce2d7
32640184
280c60b7
901c7c80
9f5cfeca
38e40067
001295dc
00412f5c
aabc12c3
00f70b47
04dc0007
0f5c0012
30c30061
22d22097
13c36026
245c1264
41471e79
24d20594
204604c3
245c0293
32c31e24
4010341c
14946207
1e69045c
10940007
90c30097
0002931c
04c30b54
41462046
0b59c0bc
fe8b101c
00f701c3
331c1eb3
09944010
30c30097
059461c7
1e69345c
ec356027
0104323c
245c69f2
46f21e71
93c36097
0001931c
2007e194
04c31654
0b3eeebc
409706d2
602732c3
000b52dc
1404345c
09547287
540c04c3
27c33900
0b514abc
d2940007
93c36097
000c931c
03c35754
218713c3
23c319b4
42546047
204710c3
000707b4
40272d54
000b24dc
00971273
208710c3
30c34a54
2b146087
216710c3
000a64dc
40970933
61e732c3
000912dc
21e712c3
32c309b4
295461a7
21c712c3
000964dc
409708f3
628732c3
12c35b54
395422c7
620732c3
0008a4dc
8f5c0e53
04c30007
25c316c3
32bc37c3
0ed30b5a
16c304c3
37c325c3
0b4c22bc
04c30df3
25c316c3
a4bc37c3
0d130b60
16c304c3
37c325c3
0b49e6bc
04c30c33
25c316c3
f6bc37c3
0b530b71
16c304c3
37c325c3
0b4c5cbc
04c30a73
25c316c3
9ebc37c3
09930b63
16c304c3
37c325c3
0b5a5ebc
00a608b3
1e6d045c
200604c3
0b3eeabc
740c06d2
1de4145c
740f6c80
1e24245c
4004323c
3e546007
6a9232c3
1e27345c
8f5c0733
40060007
04c34077
25c316c3
b2bc37c3
00f70b4f
1118301c
0000311c
680c4c0c
60076dec
686c1a15
366404c3
04c302d3
25c316c3
8cbc37c3
01d30b66
16c304c3
37c325c3
0b6f98bc
04c300f3
25c316c3
1ebc37c3
00f70b75
10c300d7
08943287
7f85740c
0093740f
fecd301c
00d760f7
c0760496
08040f56
1f36f016
60c3fc96
92c3c1c3
804ca3c3
17948007
00803f3c
af5c6037
3f3c0027
24bc00f0
00070b45
000b04dc
20372097
0027af5c
1cc306c3
3f5c29c3
0b730079
638c6810
8ba483c3
e007f04c
3f3c5894
60370080
0027af5c
00f03f3c
0b4524bc
000770c3
000924dc
501c4097
231cfe6c
d5dc481e
383c0008
4f5cffc0
32e40079
784c3334
150d435c
6097584c
684f6085
301cb84c
311c10f8
6c0c0000
60978c0c
0040033c
4426392c
65d0301c
0017311c
140f4664
0c0c784c
0007b066
2cc36854
240c19c3
133c6880
28c3ffc0
08cbb0bc
0c71784c
29c358c3
7500480c
59c37f85
57c3740f
40370a93
0027af5c
1cc306c3
34c329c3
0b7672bc
093350c3
18c3506c
501c6500
37e4feb8
700c42b4
1cc30d00
28c31b84
08cbb0bc
686c584c
686f3884
740c59c3
740f3884
606c184c
204ca006
32e421c3
2f3c2c94
60060100
fc7e323c
800c204c
1509505c
ffc0313c
20776037
143c06c3
35c30040
0b7672bc
301c50c3
311c10f8
6c0c0000
8c4c584c
392c080c
301c4426
311c65d0
46640017
2006784c
784c2c0f
00732c4f
fece501c
049605c3
0f56f876
00000804
1f36f016
50c3fe96
1404405c
431c8ad2
0754febd
feb9431c
92870454
0016c4dc
3bc0b53c
0740753c
2a00a53c
29c0953c
84c38006
0040cf3c
1e51355c
19546047
03b46047
00b369d2
23546067
33546087
fed3401c
355c2a13
341c1e24
69f24000
20a605c3
0b4e04bc
000740c3
001443dc
9f5c776c
05c30007
27c313c3
c6bc3ac3
40c30b4b
74dc0007
40660013
1e55255c
1e24355c
4000341c
05c36af2
14e3155c
0b4e04bc
000740c3
001263dc
055c0086
17b01e55
200605c3
0b3eeabc
4d540007
1e09155c
49942007
14e3655c
16c305c3
0b4900bc
000740c3
0010e3dc
17ac776c
05c36c00
23c313c3
bcbc36c3
00070b5d
000fd3dc
1e24355c
2000341c
355c6ad2
602715c9
77ac0694
15a3055c
77af6c00
15c9355c
08946047
15c1355c
04546147
610577ac
776c77af
6c0017ac
14e3255c
1501455c
0007bf5c
13c305c3
b2bc34c3
40c30b5f
23dc0007
255c000d
255c14e3
60261dc7
1e0d355c
1501355c
b2dc62a7
62a70008
628704b4
02b30694
065462c7
785462e7
fec9401c
355c17d3
341c1e24
60074000
05c37594
27c3376c
b2bc778c
0db30b77
26e605c3
0b47aabc
08d240c3
1e24355c
4000341c
52dc6007
355c000a
341c1e24
67d20010
4801255c
401c44d2
1333fe7a
200605c3
0b3eeabc
355c0ed2
6bd21e81
1de4355c
6c0017ac
155c77af
65a014e3
14e6355c
14e3355c
04546027
feab401c
255c1013
32c31e24
011c0606
30830800
111c2406
01c30800
0a9430e4
200632c3
1000111c
64f23183
fe86401c
77ac0d53
77af6025
255c4026
05c31e05
08bc2046
40c30b8b
5d940007
355c346c
341c1e24
66f20010
65a0201c
0017211c
201c00b3
211c65a4
05c30017
0b569ebc
05c300d3
27c3376c
0b5a7ebc
800740c3
08331a54
178c776c
05c30037
27c313c3
60bc3cc3
40c30b49
33540047
33740007
67f26057
fea9301c
1407355c
057343c3
27546667
155c2006
d7ac1e55
32c3578c
031463e4
03f38006
582008c3
14e3355c
103423e4
255c4086
05c31e55
eabc2006
00070b3e
ffeb22dc
1de4055c
77af7820
2006d593
1e55155c
401cd513
0073fec8
fec7401c
029604c3
0f56f876
00000804
0336f016
61c340c3
93c382c3
680c41d7
6047e006
60060454
e026640f
1404345c
febd331c
72870354
60060494
1407345c
1404045c
031c04d2
5694feb9
1e79345c
27546147
c4bc04c3
00270ba3
345c2254
72871404
1fc64994
04c308f3
0b787ebc
1407045c
15150007
fea9031c
031c3c54
3a94fecc
1e24345c
8000201c
0001211c
60073283
301c3154
345cfe73
05731407
0544545c
e254a007
051585e4
61d74026
58c34c0f
145c180c
03f20524
0093380f
b0bc25c3
39c308cb
345c6bf2
6ea00544
0547345c
0524345c
345c6e80
ebf20527
0544345c
245c68f2
45d203e1
17c304c3
0b4e4abc
c07605c3
08040f56
fe967016
940ca197
c037c1d7
c077c0cc
12c301c3
34c323c3
0b1c86bc
03f40007
0006140f
0e560296
00000804
3f36f016
60c3f496
02f70006
165c2006
365c1ea5
610715d9
60061094
73c36177
15f9465c
b4dc8007
365c0053
6c0c0764
69946007
00052d9c
0a546047
63546107
41774006
a2c372c3
db9c52c3
365c0004
60070644
005162dc
0684365c
12dc6007
365c0051
600706c4
301c1794
311c10f8
6c0c0000
0664265c
023c8c0c
392c0020
301c41e6
311c62f0
46640017
06c7065c
22dc0007
365c0050
60070704
301c1794
311c10f8
6c0c0000
0664265c
023c8c0c
392c0020
301c41e6
311c62f0
46640017
0707065c
82dc0007
265c004e
465c0644
565c0664
365c0684
603706a4
0704065c
363c0077
60b70e40
06c4165c
363c20f7
61370dc0
12c306c3
35c324c3
0b6ceabc
06930177
1fc4365c
1d946007
10f8301c
0000311c
8c0c6c0c
392c0a06
301c44a6
311c62f0
46640017
1fc7065c
42dc0007
392c004b
4764265c
0ace5ebc
00070177
004ad4dc
2021265c
61776006
12944007
165c06c3
16bc1fc4
01770b6d
128704d2
0049d4dc
065c0026
21572025
64dc2007
40260049
1ea5265c
15d9365c
e2dc6047
6107001a
003394dc
0100101c
801c22f7
811c10f8
28c30000
8c0c680c
392c01c3
301c44c6
311c62f0
46640017
0007a0c3
004732dc
1fc4065c
2f3c1ac3
4cbc02c0
50c30ad1
fe9e401c
e0068177
74dc0007
9f5c0045
365c0164
602715e1
60670554
004084dc
a2b707d3
680c28c3
001c8c0c
392c0098
301c4146
311c62f0
46640017
0007198f
004392dc
79af6146
265c392c
e6bc4764
01770b0e
04dc0007
365c0043
0c0c0764
02801f3c
6c4c598c
0abeb4bc
00070177
004234dc
4cbc198c
00070b1c
01770515
1b9c75c3
365c0004
c0c31ed2
fe67101c
e0062177
13dcc3e4
07730041
48c3a2b7
8c0c700c
392c0a06
301c44a6
311c62f0
46640017
0007198f
003fd2dc
39af24a6
265c392c
5ebc4764
01770ace
44dc0007
365c003f
0c0c0764
02801f3c
6c4c598c
0ab1a4bc
00070177
003e74dc
78bc198c
40c30ace
72bc198c
20c30ace
1ee2365c
001cc4c3
0177fe66
23e4e006
003d63dc
0040393c
393c6237
b3c30060
06c3bc84
0b3ed2bc
b21c03d2
1b3c0002
21b70090
88bc06c3
01770b4d
e4dc0007
365c003b
83c30444
0464265c
80668284
8d2d38c3
00a10f5c
065c0d4d
b0bc1fc4
18c30b4a
2f5c056d
458d0161
00d0083c
42d71ac3
08cbb0bc
943c82d7
06c300d0
0b3ed2bc
0007782c
235c2254
08c30a89
40a119c3
782c81c5
0a91135c
782c2221
0a89335c
0f546087
05b46087
14dc6047
01730034
055460a7
b4dc60c7
6e330033
6e13a0c6
6dd3a0a6
6d93a086
0a91335c
6027a086
a1060294
32c34217
23c36805
d01c61f7
d11c10f8
4dc30000
8c0c700c
392c02c3
301c44c6
311c62f0
46640017
000770c3
003562dc
133c784c
44060100
08cbb0bc
073c784c
133c0200
44060300
08cbb0bc
0400073c
0090183c
b0bc4217
05c308cb
0b23f0bc
0587065c
640c1dc3
392c8c0c
301c44c6
311c62f0
46640017
065c30c3
00070567
0032c2dc
0584265c
05c34037
41d717c3
0b257cbc
00070177
003264dc
365c99d1
602715e1
001ec4dc
d2bc06c3
00070b3e
0dc34154
8c0c600c
0200001c
44c6392c
62f0301c
0017311c
50c34664
52dc0007
782c0030
0a89235c
019e301c
10544087
05b44087
40476b06
01530a94
019f301c
065440a7
01a0301c
025440c7
05c36006
0564165c
0584265c
0ab594bc
0587065c
10f8301c
0000311c
8c4c6c0c
0564065c
44c6392c
62f0301c
0017311c
565c4664
1b8b0567
198418c3
0b3f08bc
0002921c
365c33d3
465c0664
6e0006a4
065c60c5
6c0006e4
565c6277
20061e24
4000111c
b3c35183
0000c01c
4d94a007
301ca2b7
311c10f8
6c0c0000
001c8c0c
392c0098
301c4146
311c62f0
46640017
0007198f
002b72dc
59af4146
265c392c
e6bc4764
01770b0e
e4dc0007
365c002a
0c0c0764
22dc0007
1f3c002a
598c0280
b4bc6c4c
01770abe
e4dc0007
198c0029
0b1c4cbc
04150007
75c30177
365c52d3
101c1ed2
2177fe67
03e475c3
0028e3dc
8257c0c3
604534c3
b084b3c3
d2bc06c3
03d20b3e
0002b21c
00902b3c
41b712c3
88bc06c3
01770b4d
64dc0007
365c0027
83c30444
0464465c
08c38484
41861bc3
4abc36c3
065c0b44
183c0663
08bc0090
083c0b3f
165c00b0
265c0644
b0bc0664
465c08cb
343c0664
065c00b0
28c306a3
08bc2980
81a50b3f
0e0038c3
0684165c
06a4265c
08cbb0bc
06a4065c
065c9000
28c306e3
08bc2a00
80450b3f
0e0038c3
06c4165c
06e4265c
08cbb0bc
065c94c3
908406e4
1e24365c
111c2006
31834000
e15763d2
06c31c93
0b3ed2bc
0007782c
035c2754
28c30a89
0a2149c3
0010493c
135c782c
2a210a91
335c782c
60870a89
60871354
604704b4
02130994
045460a7
049460c7
a0c63e13
201c3df3
4177ff7b
a7c3e006
a0a63613
a0863cf3
335c3cb3
a0860a91
02946027
0cc3a106
198418c3
0b3f08bc
a3c36257
0040a21c
10f8d01c
0000d11c
700c4dc3
0ac38c0c
44c6392c
62f0301c
0017311c
70c34664
32dc0007
784c001d
0100133c
b0bc4406
784c08cb
0200073c
0300133c
b0bc4406
073c08cb
183c0400
42570090
08cbb0bc
f0bc05c3
065c0b23
1dc30587
8c0c640c
44c6392c
62f0301c
0017311c
30c34664
0567065c
92dc0007
265c001a
40370584
17c305c3
7cbc2ac3
01770b25
74dc0007
921c001a
99d10002
335c782c
a0c30a91
59946027
d2bc06c3
a0c30b3e
53540007
600c0dc3
001c8c0c
392c0200
301c44c6
311c62f0
46640017
000750c3
0017e2dc
235c782c
301c0a89
4087019e
40871054
6b0605b4
0a944047
301c0153
40a7019f
301c0654
40c701a0
60060254
165c05c3
265c0564
94bc0584
065c0ab5
301c0587
311c10f8
6c0c0000
065c8c4c
392c0564
301c44c6
311c62f0
46640017
0567565c
0000a01c
e0060213
415757c3
14dc4007
61570011
83c361b7
c3c393c3
73c3b3c3
0073a7c3
81778006
065c0046
365c1ea5
604715d9
61073254
365c5494
602715e1
60670454
02534e94
0764265c
0564165c
0584465c
0380363c
798c6037
080c6077
684c00b7
000660f7
265c0693
465c0564
593c0584
363c0020
60370380
0077198c
20b72006
213720f7
12c306c3
48c324c3
40bc7280
04930b6d
335c782c
60270a91
065c2094
20061e24
4000111c
00070183
265c1894
165c0764
465c0564
363c0584
60370380
6077798c
60b7680c
60f7684c
06c30137
38c324c3
74bc3984
01770b7a
0157a006
54dc0007
20660009
1ea5165c
15d9365c
1a546047
4e946107
15e1365c
21546027
ff7b201c
a0064177
14dc6067
1b8b0008
198418c3
0b3f08bc
3ca479cc
8197b384
81b79180
782c06f3
0a91335c
32946027
1e24365c
111c2006
31834000
2a946007
10f8301c
0000311c
8c0c6c0c
392c19cc
301c44c6
311c62f0
46640017
000750c3
18c35454
59cc1984
08cbb0bc
465c79cc
065c0564
00370584
2077398c
15c306c3
34c323c3
0b71bcbc
41570177
3f944007
a0060053
365c6086
365c1ea5
60c715d9
61070354
201c0d94
4177feb8
600738c3
08c32e54
41861bc3
4abc36c3
06c30b44
419718c3
04bc6006
01770b50
1f940007
465c80a6
365c1ea5
01970464
365c6c00
365c0467
341c1e44
65f20008
d6bc06c3
01770b44
165c2086
01331e6d
ff7b301c
e0066177
007357c3
81779066
0fd20ac3
10f8301c
0000311c
8c4c6c0c
392c0ac3
301c44c6
311c62f0
46640017
301cefd2
311c10f8
6c0c0000
07c38c4c
44c6392c
62f0301c
0017311c
a0074664
301c3054
311c10f8
6c0c0000
05c38c4c
44c6392c
62f0301c
0017311c
04334664
943ca0e6
93330010
943ca0e6
c4130010
21773066
50660093
e0064177
f873a006
fec1401c
013334c3
01771066
201c0113
4177fec3
70660073
e0066177
f833a006
7ebc06c3
01570b51
fc760c96
08040f56
0f36f016
70c3f996
21b72006
205c4006
305c1ea5
341c1e24
51c30003
82dc6047
20260024
0b3eeabc
0400101c
101c03d2
07c30466
0b4d88bc
000760c3
