854ca4ec
7009444c
3b946027
0361355c
37946007
ca8c70cc
30e406c3
10ab32b4
080c303c
6d0057cc
7069708f
12946027
323c50cb
03e4080c
323c0df4
17cc100c
70ef6c00
0379255c
40f74072
00613f5c
70cb01d3
d7cc6112
70ef6f00
0379055c
241c20c3
40b700fe
00413f5c
037d355c
d04dc006
6e0c660c
204607c3
d00d3664
708c57cc
423432e4
0361655c
3e94c007
60277009
10cb3b54
080c103c
70ef6500
0053845c
080c383c
6d0057cc
7069708f
17946027
15f481e4
100c303c
6c0017cc
155c70ef
20720379
2f5c2077
255c0021
07c3037d
211230cb
09874abc
02f306c3
611270cb
6f00d7cc
055c70ef
10c30379
00fe141c
2f5c2037
255c0001
07c3037d
4abc30cb
00060987
00260053
80760496
08040f56
0736f016
50c3fd96
40772364
60373364
0430e04c
28c32450
40576949
0487623c
03a0a83c
4e946047
375c6026
602c0185
6c2c6f00
4d4d4026
6f00602c
29c36c4c
0243225c
0246235c
6f00602c
40266c2c
602c4ccd
0c2c6f00
82bc18c3
74ac0942
4c0d4026
400674ec
0395235c
235c74ec
3f5c039d
7e2d0021
6f00742c
6b0c4c4c
6b0f6c72
6f00742c
29c36c4c
4f6d4b69
6f00742c
28c36c2c
0279225c
027d235c
6f00742c
033c6c2c
1ac303a0
097fb6bc
6f00742c
28c36c2c
0333225c
0336235c
60ec08f3
235c4006
60170395
0487433c
6e00602c
40466c2c
3f5c4d4d
60b70001
6e00602c
2f5c6c4c
4cad0041
00413f5c
602c7e2d
6c2c6e00
4ccd4026
4e00602c
082c6f00
82bc2c2c
60060942
0185375c
402674ac
742c4c0d
4c4c6e00
6c726b0c
742c6b0f
6c4c6e00
4b6929c3
742c4f6d
6c2c6e00
225c28c3
235c0279
742c027d
6c2c6e00
03a0033c
b6bc1ac3
0396097f
0f56e076
00000804
0f36f016
a0c3fa96
0070c00c
b84c78b0
3970f98c
313c3629
582c0487
6c2c6d00
568c6d49
60946027
0026323c
084b133c
2f5c2037
560d0001
60257d0c
7c497d0f
4b356407
88092bc3
84f27a0c
20c66e0c
6eac0c13
36643629
355c6006
36290135
0487313c
6d00582c
6b0c4c4c
6b0f6c92
6c293bc3
1f5c6137
362d0081
323c4117
382c0487
6c2c6c80
4d4d4046
39c32006
15712c2d
486928c3
01e5255c
646918c3
400677ee
255c560d
255c0185
02c301cd
094a24bc
033c788c
155c22a0
255c01e1
febc01f1
7a0c097b
0ac36e0c
36642166
3bc32006
0cb32c0d
0010133c
2f5c20f7
5c4d0061
123c0bd3
20b70024
402624d2
0093560d
00413f5c
19c3760d
64076429
3bc34935
7a0c8c09
6e0c87f2
20a60ac3
04c33664
6eac08f3
36290ac3
1bc33664
21772429
00a12f5c
313c562d
582c0487
4c4c6d00
6c926b0c
60066b0f
0135355c
36297c4d
0487313c
6d00582c
60268c2c
956f714d
155c3069
706901e5
402677ee
0185255c
01cd255c
24bc02c3
043c094a
155c05e0
255c01e1
febc01f1
7a0c097b
0ac36e0c
36642166
3bc32006
00262c0d
133c0133
20770010
00213f5c
682d29c3
06960006
0f56f076
00000804
0136f016
80c3f896
136472c3
a00c2177
d4cc94ec
41374809
4c544047
32c34117
05b46047
40274dd2
04d30994
32c34117
59546067
608732c3
00266b54
950c0ef3
70cd7ca9
00812f5c
69d250ed
698c28c3
1f3c6c0c
366401c0
708f61d7
000c375c
70af6112
10cf0006
41725989
3f5c40f7
798d0061
356c0b73
044d1d29
323c4157
142c0487
3f5c4c00
61b700a1
0f5c684c
0cad00c1
00c13f5c
682c646d
133c03c3
00bc05e0
19890942
00b70372
00412f5c
615705b3
0487433c
6e00742c
40066c2c
760c4ced
12c36e0c
760c3664
08c36eac
00a12f5c
366412c3
6e00742c
00066c2c
04730ccd
bebc15c3
345c097e
60270361
760c0694
08c36e0c
36642006
03c37989
00fd041c
2f5c0077
598d0021
798901d3
241c23c3
403700f7
00013f5c
760c798d
41576e8c
366412c3
08960006
0f568076
00000804
fe96f016
136470c3
c00c2077
0487313c
ad00582c
6e0c7a0c
36642006
46ec344c
000632c3
0004011c
60073083
32c31054
66ef7292
8e6c7a0c
2f5c07c3
12c30021
60264046
744c4664
02730046
000632c3
0008011c
6ed23083
739232c3
07c366ef
00212f5c
404612c3
09a7d2bc
0026744c
744c0d6d
32c34d69
60377fe5
00013f5c
08b46027
6eac7a0c
2f5c07c3
12c30021
02963664
08040f56
0136f016
60c3fa96
600c81c3
8d0cac4c
3089ee0c
20272137
70a92b94
22356047
0119255c
400740f7
3f5c1d94
70ad0061
00611f5c
12c3308d
00813f5c
76bc23c3
700c0941
21772117
37546007
00812f5c
01e5235c
06c37e2c
3664300c
700f60d7
233c00f3
40b70010
00413f5c
350c70ad
211c4006
1283ffff
20072077
70891694
13546027
133c768c
20370024
402628d2
3f5c560d
355c0021
00f30135
00011f5c
4026360d
0135255c
01c9055c
094a6abc
0c0f38c3
21772006
00a12f5c
069602c3
0f568076
00000804
ff967016
a00c61c3
00403f3c
233c4006
560cfe7e
1fc3892c
36c34046
14cc4664
36bc2017
01960943
08040e56
ff967016
a00c61c3
00403f3c
233c4006
560cfe7e
1fc3892c
36c34086
14cc4664
36bc2017
01960943
08040e56
ff963016
3f3ca00c
40060040
fe7e233c
892c560c
40661fc3
46646006
201714cc
094336bc
0c560196
00000804
fe963016
80ac51c3
303c04eb
607700f4
00212f5c
6469514d
4026700d
203c440d
40370304
602644d2
0093710d
00012f5c
02bc510d
10ee0984
70ce750b
0c560296
00000804
ff96f016
72c340c3
636461c3
6c0c618c
36641fc3
d68ea017
6c6b70cc
6c802017
6017744f
0130233c
8c6b70cc
75af6a00
0100363c
2006744e
400636ae
75ac0193
8d218226
0010323c
236423c3
fff0363c
636463c3
0026d5f2
384b203c
0014103c
0067323c
60456c80
453c8006
323c371d
6c800037
20066045
3b9d153c
00c70025
07c3ec94
e0bc15c3
01960942
08040f56
0304303c
008e001c
001c6bd2
66070097
001c0754
64070091
001c0394
08040099
326430c3
00ae001c
0c5460a7
085460c7
008e001c
065460e7
61070006
001c0394
08040096
313cfe96
6037ff60
00013f5c
07b46047
333c628c
6672304b
01336077
4c69600c
341c32c3
233c001f
40770605
00213f5c
029603c3
00000804
ff963016
23641364
4f5c3264
60270081
42274994
313c05b4
60070084
46c74894
313c0ab4
67f20024
0099501c
4086a00e
0fd34037
09b44a67
0044313c
501c66f2
a00e0097
feb34106
70358047
016f231c
313c07b4
64f21004
0099201c
231c07d3
07b40228
2004313c
201c64f2
08130097
5c358087
02a7231c
31c308b4
1000341c
0099501c
42546007
03fd231c
31c34fb4
2000341c
4a946007
0097501c
41e6a00e
4227f913
313c09b4
66d20084
0096501c
4066a00e
4367f7d3
313c07b4
501c0104
6007008e
8047b494
4f273135
313c09b4
66d24004
0096201c
6146400e
231c04b3
09b400b7
8004313c
201c66d2
400e008e
03536166
1a358087
00e0231c
31c30ab4
4000341c
501c66d2
a00e0096
f23341c6
0153231c
31c30bb4
60073164
201c0715
400e008e
603761e6
a0060073
2f5ca037
02c30001
0c560196
00000804
ff963016
426440c3
23641264
026403c3
fff0503c
3f5ca037
60270001
202755b4
81072a94
81670554
81e70354
323c0594
6312ffe0
80870233
81470554
81c70354
323c0594
6212ffe0
80e70273
81a70354
323c0894
333c180c
333c02b7
013381cb
045480c7
81876006
323c0494
3364100c
02536265
03548147
079481c7
ffe0323c
333c6212
01130037
03548167
079481e7
ffe0323c
03c36312
06f30364
05948087
fff0323c
04736312
035480e7
049481a7
180c323c
8187fe33
323c2794
333c100c
61450037
00070293
80a71f94
323c0494
01b3480c
079480c7
100c323c
0037333c
00b36045
069480e7
180c323c
036403c3
81070253
323c0994
6212ff60
0037333c
00b4321c
0006fe93
05948067
fff0323c
00b36212
08948047
100c323c
0037333c
036403c3
802700b3
001c03b4
008500ca
0c560196
00000804
fe967016
61c350c3
226443c3
42644037
6c0c618c
00401f3c
60573664
2f2e2026
40066c4f
01e5235c
54cc8f4e
21c32869
4d004205
00011f5c
00df123c
02c3780f
0e560296
00000804
70c3f016
608c000c
c14ca18c
135c2a46
4a66017d
0185235c
135c2926
4be6018d
0195235c
435c8846
8a86019d
01a5435c
01ad235c
235c4886
48a601b5
01bd235c
435c8ac6
135c01c5
286601cd
01d5135c
01dd235c
135c2006
41a601e5
135c4c4d
8026014d
0155435c
235c4206
43c6015d
40a64ded
2e0d4cad
235c4006
4e8d10e6
4ccd5f46
4ced4146
03fd201c
1106235c
2dcd2ead
e8c95e2c
610ceecd
616c2d0d
616c8c4d
2000201c
201c4cae
548e0200
74ae6246
348d94ed
78ce58ae
0f56386d
00000804
fd961016
026443c3
126400b7
22642077
05b44027
700d6006
17130066
40676026
40470454
60060494
13f3700d
31c32057
60377fe5
00013f5c
85dc6027
60970008
35946007
06944147
700d6026
0080001c
41c713b3
60260694
001c700d
12d300e7
04944087
700d6026
416710f3
60260694
001c700d
115300be
069441e7
700d6026
015a001c
40e71073
60060594
0466700d
41870fb3
60060594
0fa6700d
41a70ef3
60067494
001c700d
0e1300b9
31c32097
49946027
06944087
00413f5c
07a6700d
41470cb3
3f5c0794
700d0041
0176001c
41c70bb3
3f5c0794
700d0041
02ae001c
41070ab3
60260594
0b46700d
416709f3
60260694
001c700d
0913022f
069441e7
700d6026
0404001c
40c70833
60060594
0826700d
40e70773
60060594
0be6700d
418706b3
60060694
001c700d
05d3016d
069441a7
700d6006
0221001c
200604f3
0473300d
700d6006
20570413
1d942007
069440a7
00211f5c
01a6300d
40c702f3
1f5c0694
300d0021
021302e6
069440e7
00211f5c
0426300d
41070133
1f5c0694
300d0021
00530326
03960006
08040856
20c331c3
32642364
059460a7
41470006
01b30f35
059460c7
42870006
00f30935
60e70026
00060594
023543c7
08040026
326430c3
22641364
2d946027
14544067
045440a7
48944027
31c30373
2000341c
03fd001c
45546007
341c31c3
001c1000
600702a7
313c3e54
001c2004
60070228
313c3854
001c1004
6007016f
313c3254
0a660044
2d546007
0024313c
600706c6
04f32394
13544067
045440a7
20944027
31c302f3
001c3164
60070153
31c31a74
4000341c
00e0001c
13946007
8004313c
00b7001c
313c6ef2
0f264004
313c6af2
03660104
313c66f2
02260084
000662f2
00000804
698c400c
20062cef
2ccd2d0f
6c0c684c
2cad2206
6e0c6a0c
366420c6
00000804
40c31016
414c000c
200628af
68ab290f
07ff331c
301c0535
686e03ff
2fe60073
6006286e
684d682d
6c0c604c
2cad2206
6e0c620c
204604c3
08563664
00000804
31c3fe96
60773264
40372264
2057604c
202724d2
02131594
00011f5c
40172e2d
202712c3
2f5c0594
4ccd0001
1f5c0133
2ccd0021
60ac00b3
00012f5c
02964c2d
00000804
0136f016
50c3fa96
82c361c3
004ce0ec
175c800c
21c30361
40375fe5
00013f5c
07b46047
8b33201c
009e211c
0173506f
282b416c
341c31c3
70120fff
280b706f
706f31a3
21c3306c
301c2364
311c0284
4c0e4107
808c213c
4c0e6045
308f228c
0361375c
295460a7
0ab460a7
20546047
72b46047
70546007
09946027
61270153
60e704b4
09b36934
52356187
04f34026
4d0c750c
341c6520
23063fff
331c2077
03351fff
60776106
00211f5c
600602d3
754c702d
06f34c49
4049156c
11944007
652040cc
003f341c
20b72306
033563e7
60b76106
00411f5c
4006304d
07d34177
0f944027
652040cc
1fff341c
20f72306
0fff331c
61060335
1f5c60f7
fdb30061
2a944047
652040cc
3fff341c
21372306
1fff331c
61060335
1f5c6137
fbb30081
4cc9758c
440d18c3
61776006
784c02f3
60276f69
582c1194
03a0323c
32c3704f
213e133c
241c21c3
4c0e7fff
235c782c
502d0279
2006fd53
2f5c2177
02c300a1
80760696
08040f56
00870364
01071654
01671454
01471254
01e71054
01c70e54
303c0c54
233c0036
303cfff0
7fe50096
033c32a3
0053f88c
08040026
630d6006
636d632d
634d638d
62cd62ad
01c5305c
0804628d
0736f016
40c3f996
2177200c
2450a48c
6c0c618c
01801f3c
c1973664
c86f29c3
7aae6006
6c6b70cc
6c802197
733c784f
f9af0100
0140a33c
153c0ac3
56691270
08cbb0bc
823c5669
b6290040
a157a137
093c760c
21170420
a0a629d2
00055f5c
101c8ecc
60064408
20a60153
00051f5c
101c8ecc
5f5c8818
35c30081
30c34664
233c3264
40f7180c
00615f5c
2006bc0d
533c3c2d
a0b7ffd0
00413f5c
ffc0283c
12b46027
180c323c
60776172
00213f5c
073c7c4d
1ac30030
08cbb0bc
fff0383c
836483c3
323c00b3
6172180c
383c7c2e
784e0100
386f2006
686c29c3
0146835c
e0760796
08040f56
0336f016
72c360c3
800c1364
105050ec
76c958c3
a4dc6027
20470008
720c0b94
20066eec
522c3664
6025690c
0006690f
325c1093
60270361
20676d94
21470b54
21c70954
20870754
21670554
21e70354
722c6194
40254d2c
110c4d2f
6ef26089
0026800c
69948007
6c6c798c
17c306c3
58c33664
04c3942f
313c0c13
3364ffd0
35e4a026
a0460235
78cc000c
204c4c69
133c6880
7c4c0100
923c4980
7c0b0130
5f6523c3
0580600b
2e8039c3
b0bc4aa0
710c08cb
080b4c0c
60803c0b
6ea07f65
710c680e
08cb4c0c
60803c0b
6ea07f65
798c68ce
06c36c6c
366417c3
28c36006
710c682f
a0064c0c
0026ac0f
01e5025c
6e2c720c
12c306c3
710c3664
2cad2006
2c8d710c
200606c3
76bc4026
05c30941
b6bc0293
798c0948
06c36c6c
366417c3
28c36006
03c3682f
618c0113
17c36c6c
00063664
142f58c3
0f56c076
00000804
0136f016
60c3ff96
1cb0e00c
bc4c9cec
0119355c
233c68d2
4037fff0
00013f5c
011d355c
0948b6bc
0361445c
3e5480c7
06b480c7
09548047
7b9480a7
80e70313
81676a54
0d937694
202606c3
76bc4006
7d4c0941
2c8e2006
20e606c3
76bc4026
7e0c0941
06c36e0c
0c532066
566c740c
06c34caf
40062066
094176bc
6e0c7e0c
20e606c3
740c3664
21c32cac
301c2364
311c0288
4c0e4107
808c213c
4c0e6045
69cc5e2c
69cf6025
06c30893
40062046
094176bc
20067d8c
06c32cce
402614c3
094176bc
6e0c7e0c
210606c3
7d8c3664
01c9055c
46f24cc9
6abc940c
10af094a
6abc0113
740c094a
4c124ca9
4caf4100
2cac740c
236421c3
0288301c
4107311c
213c4c0e
6045808c
5e2c4c0e
60256a2c
01f36a2f
6a0c5e2c
6a0f6025
18c300b3
60276409
7e0c0694
06c36e0c
36642146
80760196
08040f56
1f36f016
90c3fa96
21371364
5450a00c
04301ac3
6abc0006
28c3094a
233c684c
19c30130
2c6964cc
375ce880
233c0074
303c188c
69a0108c
7fff341c
28c37d4e
31c3280b
680e6045
335c74ec
61770361
3b946027
d6bc950c
075c0949
18c300b7
32c3440b
640e6085
73c37c6b
0400741c
e007e0f7
762c1254
40254d4c
1f5c4d4f
308d00a1
200609c3
76bc21c3
10110941
2ac36006
18f3682f
00611f5c
3f5c308d
28c300a1
01e5325c
6e2c760c
18c309c3
40d73664
442f1ac3
12c309c3
00a13f5c
76bc23c3
15f30941
21c32157
09544127
04dc2167
74ac000a
60276c09
0009b4dc
3ac32006
012d135c
6a6c562c
6a6f6025
23c37d0b
1fff241c
143c47c3
31c3073e
fff8341c
c23c6152
411779ac
0487623c
6f00742c
27c30c2c
62327c4b
033e123c
71ac313c
b0c3600e
680b17c3
241c23c3
323c03ff
213c110c
323c043e
b21c41ac
2bc30002
27c3680e
6832640b
053e123c
41ac313c
1f5c604e
3ac30081
742c2e2d
6c4c6f00
41c33009
0007441c
1f5c80b7
2cad0041
6f00742c
480b6c2c
40774832
00212f5c
742c4d6d
6c2c6f00
2cce3ccb
6f00742c
6c4c8c2c
cc18201c
0206235c
6f00742c
20266c2c
74ac2ccd
60376c09
0b946027
6f00742c
8f716c4c
1f5c74ec
135c0001
0173039d
4026758c
3ac34c2d
01c9035c
20721cc3
094aa8bc
1ac34006
012d215c
440b1bc3
341c32c3
42660080
458662f2
3c0c34c3
2f7e133c
2c2f3c2c
0323145c
341c31c3
323c03ff
345c51ac
29c30326
6c6c698c
18c309c3
20063664
2c2f3ac3
f8760696
08040f56
0736f016
50c3fe96
5a10c00c
18b038f0
706c984c
68d273c3
2c096dac
341c31c3
733c0078
b6bc188c
7abc0948
30c30949
60273264
345c5854
68d20111
fff0233c
3f5c4037
345c0001
306c0115
12542007
325c29c3
61670361
28c30794
60276809
e0470994
758c0794
05c36c4c
20063664
29c3306f
0361325c
15546087
04b46087
28356047
61670113
61671954
61872314
04132a94
202605c3
76bc21c3
1ac30941
0113660c
202605c3
76bc21c3
2ac30941
05c36a0c
36642046
322901b3
0487313c
6d00582c
6d496c2c
04946047
245c4006
7a2c01dd
0404235c
235c4025
60060407
00736077
20772026
00212f5c
029602c3
0f56e076
00000804
fe96f016
20771264
40372264
f5248e24
00212f5c
6abc02c3
60c3094a
00013f5c
6abc03c3
70c3094a
00212f5c
96bc02c3
50c3094a
3f5c5364
03c30001
094a96bc
343c0364
62d24004
363cf324
65f20024
4e20353c
536453c3
0014363c
353c65f2
53c32710
373c5364
65f20024
4e20303c
036403c3
0014373c
303c65f2
03c32710
05e40364
201c0635
750009c4
536453c3
033c7420
0296088c
08040f56
3f36f016
b0c3fe96
426441c3
d264d2c3
29c32010
403748ec
4c9039c3
ec4c8cb0
6c0c618c
00401f3c
8f5c3664
1c710024
60cc0bc3
20576c6b
28c36c80
0486684f
633c084e
c9af0100
2a8e2286
6aae6006
305c0017
60670361
00060994
094a6abc
0020503c
0000d01c
2cc30453
60276809
80471b94
00061994
094a6abc
000650c3
094a96bc
436440c3
01c9075c
094a84bc
04e40364
353c0c35
60670034
60270354
a0250694
7eac0093
0020533c
fffc001c
0fff011c
101c5083
380e0290
68092cc3
04946027
29053d3c
7ac3780e
1153775c
0ac3f82e
1163005c
36c3184e
415c1ac3
24c31173
0003241c
036e233c
1c6c7bc3
213c200b
4c0e112c
602926c3
e0496632
11ac473c
336434c3
046e323c
175ce017
20670361
1ac30e94
22d22649
680e6a72
718c49c3
17c3e80b
373cece9
011360ac
079420e7
7d6c79c3
313c2c49
680e622c
34c3880b
8000401c
680e34a3
001b705c
36c3f8ae
233c40a9
0ac3066e
0149105c
203c01c3
4c0e412c
26ab1ac3
2cc338ee
60276809
3d3c0354
790e0074
733c36c3
253c083e
4c0e0bac
788c353c
2006792e
206f08c3
fc760296
08040f56
50c33016
842c01c3
640c8bd2
083532e4
0942f2bc
6c4c758c
14c305c3
0c563664
00000804
fd963016
819752c3
12640264
00c72037
00c72654
00470eb4
00471f54
00b707b4
35540007
12940027
00870273
03931135
08b40127
022a321c
40b74006
34340107
01670273
01871635
20262d54
321c06b3
40060222
321c0193
00730222
022a321c
20b72026
343c0433
402605e0
039340b7
321c5149
2006022a
404720b7
343c1554
200605e0
402720b7
01d30d94
00412f5c
3f5c02c3
13c30001
d6bc25c3
2006094a
60060173
03c360b7
01e1155c
01f1255c
097bfebc
2077fd93
00212f5c
039602c3
08040c56
2264fe96
0014313c
60096fd2
23c347d2
40774072
00213f5c
23c300d3
40374092
00013f5c
0006600d
08040296
40c33016
612c51c3
32c34c09
0001341c
6cd223c3
6c0c618c
740c3664
286b50cc
4c4f4c80
2c6f2006
02c34285
08040c56
22641016
8c09612c
341c34c3
6ad20001
223c600c
0c2c0487
033c6800
e0bc02c0
08560942
00000804
40c33016
602c52c3
01a0033c
b0bc4106
702c08cb
32c34f89
0004341c
746c6cf2
32c34d09
0004341c
708c66d2
4cad4086
4ced708c
08040c56
326431c3
013e201c
4107211c
00ff101c
201c280e
211c013c
680e4107
0168301c
4107311c
0006600f
00000804
301c200b
311c020e
2c0e4107
6045202b
204b2c0e
2c0e6045
6045206b
208b2c0e
2c0e6045
604520ab
20cb2c0e
2c0e6045
604540eb
08044c0e
301c200b
311c0204
2c0e4107
6045202b
404b2c0e
4c0e6045
00000804
43c33016
0264a0d7
0bf21264
680b24f2
680e6072
301c500b
311c009e
05f34107
0e940027
680b24f2
680e6172
6472680b
500b680e
00a2301c
4107311c
00470413
24f20e94
6272680b
680b680e
680e6572
301c500b
311c00a6
02334107
13940067
680b24f2
680e6372
31c3280b
0030351c
500b680e
00bc301c
4107311c
540b4c0e
4c0e6045
08040c56
0336f016
70c3fd96
61c37264
60066364
00563f5c
00463f5c
00363f5c
ac4c680c
2c5069ec
9886301c
4103311c
83c36c0b
355c8364
65f20189
2f5c4806
00930056
3f5c6806
355c0046
60270129
3f5c0794
62720053
00563f5c
3f5c00d3
62720043
00463f5c
01c9255c
0181155c
00803f3c
02c36037
00602f3c
00a03f3c
098dd6bc
00332f5c
311c6006
4c0e4107
0131255c
07944027
311c6186
4c0e4107
011342c3
009c301c
4107311c
4c0e4026
355c8006
60270139
393c0594
62d20014
e0478e72
cd720c94
c00f201c
363c4283
333c3ff4
43c3222c
00f34364
cc72e3f2
e0270093
ce720294
60277669
cb720294
311c6146
cc0e4107
0141255c
341c32c3
5006007f
38a38283
9886201c
4103211c
701c680e
711c0200
7c0b4107
641c63c3
355cf000
602701d1
355c1c94
600701a9
368c1894
236421c3
020a301c
4107311c
213c4c0e
6045808c
156c4c0e
098dc8bc
acbc164c
363c098d
7c0e0035
01138372
437226c3
0200301c
4107311c
301c4c0e
311c9880
8c0e4103
c0760396
08040f56
50c37016
026401c3
00834f5c
013e101c
4107111c
00ff601c
101cc40e
111c013c
040e4107
840e2085
542f740f
08040e56
21c330c3
22643264
009e101c
4107111c
101c6ed2
111c00a2
60274107
101c0854
111c00a6
60474107
22c50254
0010323c
33646a12
0804640e
226420c3
013e301c
4107311c
00ff001c
301c0c0e
311c013c
4c0e4107
0168201c
4107211c
341c680b
7f0507ff
136413c3
341c680b
31e407ff
63c6fcd4
4107311c
041c0c0b
08040004
41c31016
126412c3
60277249
60892494
241c23c3
313c000f
323c780c
23c359ac
301c2364
311c011a
4c0e4107
01b1245c
301c4ad2
311c010c
4c0b4107
41722364
01334c0e
010c201c
4107211c
341c680b
680efffd
08040856
fc967016
22641264
23c340b7
62172264
0604533c
a3d245c3
0200401c
375420c7
0ab420c7
2cb42087
27342067
0e542027
09942047
21270253
210704b4
06b33d34
3d352187
80f78a26
c0e612f3
a007c00d
20895354
0a1341a3
23c46097
f88c323c
0020133c
2f5c2037
400d0001
4454a007
433c60a9
0813d95b
c00dc106
208607b3
a007200d
40893954
06d342a3
65f26097
00416f5c
0073c00d
200d2026
2c54a007
423c40a9
0513d95b
600d60a6
2454a007
46a3c089
20c60433
03d3200d
412644f2
0353400d
600d6146
df86608c
608f3683
440b204c
028c301c
4107311c
442b4c0e
4c0e6045
6045444b
446b4c0e
4c0e6045
6045448b
60294c0e
20096112
61ac213c
60492006
02946307
21a32026
f1ff241c
0296301c
4107311c
a3d24c0e
8c0e6045
21c3208c
301c2364
311c020a
4c0e4107
808c213c
4c0e6045
0280201c
4107211c
3364680b
680e6072
0282101c
4107111c
0282201c
4107211c
341c640b
79d20001
433c680b
80f7384b
133c680b
20772a0b
00212f5c
3f5c406d
03c30061
0e560496
00000804
ff963016
41c350c3
326432c3
56bc6037
043c094c
78bc03e0
201c094c
211c010c
680b4107
60723364
7609680e
34c366f2
734e133c
01534145
10946027
133c34c3
201c75ce
211c0116
280f4107
15c303c3
00013f5c
30bc23c3
245c098f
301c00f4
311c010e
4c0f4107
0114245c
4c0f6085
0c560196
00000804
ff96f016
400c51c3
2629c88c
0487313c
6f80e82c
546c2c6c
8c0969ac
61ec4a8b
341c6c4c
6dd20002
602765a9
e4090a94
341c37c3
65d20001
0040323c
236423c3
602777c9
64460794
4107311c
ec0ee806
301c00f3
311c009a
28064107
77e92c0e
08946027
311c6446
101c4107
2c0e0080
301c0113
311c009a
701c4107
ec0e0080
20cb343c
612c233c
311c6586
4c0e4107
0213255c
311c6486
4c0e4107
60277669
61460994
4107311c
23644c0b
4c0e4b72
41460113
4107211c
341c680b
680ef7ff
6c29612c
10946027
335c60ec
60270451
64460b94
4107311c
2c0e2086
311c6346
5fe64107
255c4c0e
301c0203
311c80b2
4c0e4103
86a4201c
4103211c
3364680b
680e6372
01c9055c
094a84bc
01270364
966c1735
01c9055c
094a6abc
105440e4
311c6446
20264107
365c2c0e
641211c4
000f351c
11c7365c
40374006
60660073
7f5c6037
07c30001
0f560196
00000804
3f36f016
32379a96
226471b7
200651f7
0b3d1f5c
3f3c4006
81221570
5f5c9277
45030b39
7f5c9177
7f5c08a1
1f5c0b3d
2d210921
42074025
4f3cf194
04c31880
c4bc3217
a0260942
8f3cb4b7
8f5c1780
4f5c0087
14970a41
341c30c3
66f20001
17807f3c
18806f3c
7f3c00b3
6f3c1880
80271780
343c5c54
7137080c
08815f5c
826485c3
ffe0183c
1f5c30f7
74970861
7a056512
a888201c
0013211c
0f3cad00
9f3c1680
31c31570
06352207
fef0313c
3f5c70b7
29c30841
4c096980
288cb23c
1daca23c
0827af5c
08212f5c
2f5c52b7
4c0d0941
009f353c
69805297
3f5c7037
303c0801
313c00df
6ff70010
07e11f5c
32c34117
d89403e4
00e0983c
07c79f5c
07c12f5c
06354207
fef0123c
2f5c2f77
3f3c07a1
6d001570
45324c09
853cac09
8f5c192c
0f5c0787
0c0d0781
200627c3
15700f3c
0034313c
606763d2
71d72f94
a02753c3
80670f94
72170d94
85c3aca2
35c3a809
8f5c8303
5f5c0767
a80d0761
80270073
3f3c0d54
aca21680
a80985c3
830335c3
07478f5c
07415f5c
60a20113
680953c3
ae775303
07215f5c
6809a80d
a688501c
0013511c
71d70513
a02753c3
80670c94
72170a94
a8096ca2
6e376e80
07013f5c
0073680d
0b548027
16803f3c
a8096ca2
6df76e80
06e13f5c
0113680d
6809a0a2
adb7b580
06c15f5c
6809a80d
a788501c
0013511c
a80db5a2
40252025
a1942207
080c143c
5f5c2d77
353c06a1
6d37fff0
06811f5c
65127497
001c7c05
011ca888
8c000013
16800f3c
15708f3c
220731c3
913c0735
9f5cfef0
3f5c0667
28c30661
4c096980
288ca23c
1d2c923c
06479f5c
06412f5c
2f5c54f7
4c0d0a61
009f343c
698054d7
3f5c6c77
303c0621
313c00df
6c370010
06011f5c
32c34117
d79403e4
00f0853c
05e78f5c
05e12f5c
06354207
fef0123c
2f5c2bb7
3f3c05c1
6d001570
45324c09
543c8c09
ab77192c
05a15f5c
6006ac0d
0034233c
406743d2
0f3c0b94
01a21680
00803da2
2f5c0b37
5da10581
4f3c01b3
b1a21680
bda285c3
840345c3
05678f5c
05615f5c
6025bda1
e3946207
f337f2f7
07c3f377
203c17c3
413c049e
6a00041e
b0c332f7
053c57c3
4c00059e
17c3a5c3
051e313c
91c36112
47c34980
061e343c
c4c36112
57c34980
069e353c
d5c36112
07c34980
071e303c
13376312
17c34980
079e313c
33776212
6ab76980
05412f5c
f3b740f7
f437f3f7
47c307c3
5c0957c3
37c34112
009e133c
650073b7
123c27c3
6c80011e
27c353f7
019e123c
54376c80
031e243c
153c6d00
4c80039e
313c17c3
6212021e
498081c3
029e303c
69806112
2f5c6a77
60d70521
69806112
3f5c6a37
780d0501
488020d7
2f5c49f7
582d04e1
18c34009
68802409
4c803409
61127009
32d74980
63126409
1bc34980
62126409
19c34980
61126409
1ac34980
61126409
69b76980
04c11f5c
68095397
48092dc3
40774d00
69807c09
53176077
4d004809
73574077
69806c09
53d76037
62126809
49804017
74174037
41124c09
6d006017
2cc36037
61126809
49804017
2f5c4977
313c04a1
6980080c
3f5c6937
784d0481
28f72880
04611f5c
7c09386d
53d76312
6d004809
24093417
20096c80
33974c80
62126409
18c34980
61126409
70094980
49806112
61127409
68b76980
04411f5c
68092bc3
480952d7
40774d00
6c093cc3
60776980
48092dc3
40774d00
6c097357
60376980
680929c3
40176212
40374980
4c093ac3
60174112
60376d00
68095317
40176112
48774980
04212f5c
080c313c
68376980
04013f5c
2880788d
1f5c27f7
38ad03e1
28095397
48095417
3c096500
33d74c80
61126409
18c34980
61126409
60094980
49806112
63127009
74094980
69806212
1f5c67b7
29c303c1
2bc36809
4d004809
3ac34077
69806c09
53176077
4d004809
73574077
69806c09
52d76037
61126809
49804017
3cc34037
42124c09
6d006017
2dc36037
61126809
49804017
2f5c4777
313c03a1
6980080c
3f5c6737
78cd0381
26f72880
03611f5c
7c0938ed
53976112
6d004809
6c803009
4c803409
640933d7
49806112
64093417
49806112
640918c3
49806312
62126009
66b76980
03411f5c
68092bc3
480952d7
40774d00
6c093ac3
60776980
48092cc3
40774d00
6c093dc3
60376980
680929c3
40176112
40374980
4c097317
60174212
60376d00
68095357
40176112
46774980
03212f5c
080c313c
66376980
03013f5c
2880790d
1f5c25f7
392d02e1
61127c09
48092dc3
33176d00
6c802409
24093357
33974c80
61126409
33d74980
63126409
34174980
62126409
1cc34980
61126409
65b76980
02c11f5c
28c36009
4d004809
74094077
60776980
480929c3
40774d00
6c093ac3
60376980
61127009
69804017
72d76037
42124c09
6d006017
2bc36037
61126809
49804017
2f5c4577
313c02a1
6980080c
3f5c6537
794d0281
24f72880
02611f5c
2dc3396d
2cc32809
65004809
24093357
32d74c80
61126409
1bc34980
61126409
19c34980
63126409
1ac34980
62126409
33174980
61126409
64b76980
02411f5c
68095397
48095417
40774d00
69807c09
28c36077
4d004809
60094077
60376980
680953d7
40176112
40374980
62127009
40374980
61127409
64776980
02212f5c
080c313c
64376980
02013f5c
2880798d
1f5c23f7
39ad01e1
280929c3
48092bc3
1ac36500
4c802409
640932d7
49806112
64091cc3
49806312
64091dc3
49806212
64093317
49806112
64093357
69806112
1f5c63b7
7c0901c1
53d76212
6d004809
fc09f417
40096f80
f0096d00
14096f80
93974c00
61127009
58c34980
61127409
63776980
01a12f5c
080c313c
63376980
01817f5c
2880f9cd
0f5c22f7
19ed0161
21c33497
54b74025
84dc4127
301cffc3
311ca684
2c0c0013
94778006
15704f3c
16800f3c
0a212f5c
0100723c
3f5ce2b7
62070141
523c0654
a277fff0
01213f5c
68095180
e8096532
19ac873c
01078f5c
01013f5c
313c7537
b517009f
61f77580
00e13f5c
63a1f457
f477e025
0554e207
0a815f5c
faf3a80d
1f3c6006
233c1680
43d20034
0b944067
20c305a2
200319a2
4f5c41b7
519700c1
013389a1
f9a2a5a2
a177b780
00a12f5c
41a11197
62076025
6696e794
0f56fc76
00000804
0136f016
50c3e696
62c381c3
426443c3
05800f3c
24c312c3
0942c4bc
06407f3c
0b9480c7
05e00f3c
24c316c3
0942c4bc
16c307c3
00b34086
16c307c3
4e206206
0942c4bc
04804f3c
18c305c3
34c34006
099102bc
04c36006
05801f3c
d1a248c3
c1a226c3
240346c3
6f5c4477
c1a10221
4a0085a2
6f5c4437
c5a10201
62076025
7409ee94
9d2543c3
6f5c83f7
6f5c01e1
54290245
5ca632c3
63b73203
01c13f5c
024d3f5c
64c39449
c377dbe5
01a12f5c
02552f5c
43c37469
43037826
4f5c8337
4f5c0181
d489025d
566526c3
3f5c42f7
3f5c0161
94a90265
94e664c3
c2b76403
01416f5c
026d6f5c
32c354c9
627772a5
01214f5c
02754f5c
26c3d4e9
2603d066
2f5c4237
2f5c0101
7509027d
7d2643c3
81f74303
00e14f5c
02854f5c
26c3d529
41b75ca5
00c13f5c
028d3f5c
64c39549
64039be6
6f5cc177
6f5c00a1
55690295
782532c3
4f5c6137
4f5c0081
d589029d
d66626c3
40f72603
00612f5c
02a52f5c
43c375a9
80b794e5
00416f5c
02ad6f5c
32c355c9
320352a6
3f5c6077
3f5c0021
95e902b5
b06554c3
6f5ca037
6f5c0001
402602bd
02bc6817
1a960991
0f568076
00000804
6037ff96
4cbc6186
01960995
00000804
6037ff96
4cbc60c6
01960995
00000804
0136f016
80c3f996
73c301c3
426442c3
40b74206
2eb481e7
00c05f3c
24c305c3
0942c4bc
5a20c206
40a71600
17c307d4
0942c4bc
c0b705c3
17c303b3
c4bc40c6
343c0942
60770060
00212f5c
42c340b7
15008112
08d481e7
c4bc15c3
16000942
5a2015c3
15c30093
59a06097
0942c4bc
48c305c3
32c34097
079e243c
60373203
00013f5c
18c3700d
63574026
099102bc
32c34097
32035009
3f5c60b7
700d0041
80760796
08040f56
0136f016
70c3fa96
82c361c3
243c40c3
32c3079e
0006361c
2f5c6077
500d0021
00805f3c
40c605c3
0942c4bc
00e00f3c
40c616c3
0942c4bc
01400f3c
408616c3
0942c4bc
15c307c3
38c34026
099102bc
23c37009
0006261c
3f5c4037
700d0001
80760696
08040f56
3f36f016
60c3f996
407720b7
6d8c6037
00176c0c
01801f3c
20063664
153320f7
661260d7
09804097
303c2006
333c1a1d
4197088d
1b9d323c
22072025
4006f794
8d006197
723c31cc
0f810040
512c6d01
313cad00
213c998c
3203898c
508c213c
35803203
918c303c
398c203c
203c3203
3203188c
720f6580
00c0731c
27c30354
165cfc13
21370444
0464965c
0484865c
04a4c65c
04c4565c
04e4a65c
0504b65c
0524265c
61776197
e00641c3
27812157
201c6880
211ca9a8
4b810013
353c2d00
253c598c
3203318c
c98c253c
25803203
3b8335e3
2a8325c3
05803203
dc84d0c3
180319c3
39c31483
13033883
698c343c
118c243c
243c3203
3203b18c
6c006580
c8c3e085
731c2bc3
08540100
a5c3bac3
89c35dc3
43c394c3
4117f953
365c6d00
365c0447
6e000464
0467365c
0484365c
365c3984
365c0487
388404a4
04a7365c
04c4365c
365c3d84
365c04c7
6e8004e4
04e7365c
0504365c
365c3a84
365c0507
3b840524
0527365c
13c360d7
20f72025
32c340d7
32e44057
fff540dc
658c2017
01c36c2c
36642197
fc760796
08040f56
301c1016
311ca988
20c30013
0200133c
024f433c
0447425c
31e44085
6006fa94
600f602f
08040856
0336f016
70c3fd96
42c381c3
402c93c3
6d206806
3f5c6077
80b70021
023543e4
6f5c60b7
323c0041
1d800080
26c318c3
0942c4bc
71005c2c
03b467e7
04f37c2f
80379320
00014f5c
388c543c
673c8684
07c30080
402616c3
b6bc39c3
07c30996
25c318c3
b6bc39c3
441c0996
353c003f
06c3300c
298028c3
c4bc24c3
9c2f0942
0010353c
3c0c6612
7c0f6c80
c0760396
08040f56
099792bc
00000804
0336f016
91c360c3
402c82c3
03f4323c
66e7e046
e02602b4
6880380c
180c433c
300c573c
0080323c
20061980
b6bc5520
582c0942
30067900
443c2d0d
7a80088d
06c38c2f
0080163c
38c327c3
0996b6bc
400606c3
0444305c
088d333c
313c19c3
40252b9d
41070085
c076f694
08040f56
0136f016
60c3f096
82c371c3
5f3c43c3
15c30200
e0bc23c3
621c0997
06c300a8
440615c3
92bc34c3
06c30997
24c31fc3
0997e0bc
1fc307c3
c4bc28c3
10960942
0f568076
00000804
0136f016
60c3d696
82c371c3
0fc353c3
09977ebc
16c30fc3
35c327c3
099792bc
18c30fc3
e0bc25c3
2a960997
0f568076
00000804
0136f016
60c3f596
12c301c3
280783c3
70c30494
03b351c3
04b42807
51c370c3
4f3c0113
24c300c0
09983cbc
a40674c3
8ea06806
2a00353c
26c61980
b6bc24c3
353c0942
19802e00
24c32b86
0942b6bc
03532006
58807c80
40c30c09
0036461c
0f5c80b7
025c0041
8c091505
361c34c3
6077005c
00210f5c
1705025c
0010313c
1f5c6037
15e40001
06c3e674
09977ebc
163c06c3
48062a00
92bc38c3
463c0997
04c30a80
09977ebc
163c04c3
48062e00
92bc38c3
0b960997
0f568076
00000804
c0967016
61c350c3
612c6364
31c32c09
0001341c
600c66d2
6c0c6e0c
366416c3
10003f3c
233c4006
554c805e
05c3886c
2fc316c3
46646026
0e564096
00000804
be961016
612c1364
32c34c09
0001341c
41866037
67d24077
6c8c600c
60376e89
60776006
00212f5c
00452f5c
00013f5c
004d3f5c
8c6c614c
00802f3c
46646046
08564296
00000804
bf961016
612c1364
34c38c09
0001341c
80378186
600c67d2
88696c8c
40068e8d
3f3c4037
4f5c1040
433c0001
414c805e
23c3886c
46646026
08564196
00000804
bc967016
612c1364
34c38c09
0001341c
a0b7a026
1f546007
8c8c600c
c00634c3
a869c0f7
a007a077
6f5c1154
635c0021
a0d7017d
c02565c3
5f5cc037
a0f70001
60254025
00f8531c
2f5ced94
504d0061
60b76006
11003f3c
00414f5c
805e433c
886c414c
602623c3
44964664
08040e56
bf961016
612c1364
32c34c09
0001341c
80378026
67d223c3
6c8c600c
10d3235c
60376006
10403f3c
00014f5c
805e433c
000e235c
886c414c
606623c3
41964664
08040856
bf961016
612c1364
34c38c09
0001341c
80378026
600c69d2
425c6c8c
435c001b
400610d6
3f3c4037
4f5c1040
433c0001
414c805e
23c3886c
46646026
08564196
00000804
bf961016
612c1364
32c34c09
0001341c
80378026
66d223c3
6d6c600c
60064cab
3f3c6037
4f5c1040
433c0001
235c805e
414c000e
23c3886c
46646066
08564196
00000804
bf961016
612c1364
34c38c09
0001341c
80378026
600c6bd2
001b225c
80378246
6d6c45d2
40064cae
3f3c4037
4f5c1040
433c0001
414c805e
23c3886c
46646026
08564196
00000804
be961016
612c1364
32c34c09
0001341c
40374026
67d26077
6c8c600c
60776e09
60376006
00012f5c
00452f5c
00213f5c
004d3f5c
8c6c614c
00802f3c
46646046
08564296
00000804
bf967016
61c350c3
612c6364
31c32c09
0001341c
20372026
600c68d2
6c8c6e0c
36642869
40374006
10403f3c
00011f5c
805e133c
886c554c
16c305c3
602623c3
41964664
08040e56
bf963016
612c1364
32c34c09
0001341c
a02666f2
23c3a037
00f343c3
6d8c600c
8c8b4cab
60376006
10403f3c
00015f5c
805e533c
000e435c
001e235c
886c414c
60a623c3
41964664
08040c56
be967016
536451c3
2c09612c
341c31c3
c0260001
6007c077
600c2154
2e248d8c
325cf524
708e001b
002b225c
708b50ae
0800331c
23030ab4
633c32c4
c037f88c
00012f5c
007350ed
70ed6046
4004313c
64d26077
c006f324
3f3cc077
1f5c1080
133c0021
414c805e
15c3886c
602623c3
42964664
08040e56
bf963016
612c1364
32c34c09
0001341c
a02666f2
23c3a037
00f343c3
6d4c600c
8cab4ccb
60376006
10403f3c
00015f5c
805e533c
000e435c
001e235c
886c414c
60a623c3
41964664
08040c56
bf961016
612c1364
34c38c09
0001341c
80378026
600c6bd2
425c6d4c
8cce002b
001b425c
40068cae
3f3c4037
4f5c1040
433c0001
414c805e
23c3886c
46646026
08564196
00000804
be961016
612c1364
32c34c09
0001341c
40374026
67d26077
6c8c600c
60776d29
60376006
00012f5c
00452f5c
00213f5c
004d3f5c
8c6c614c
00802f3c
46646046
08564296
00000804
bf961016
612c1364
34c38c09
0001341c
80378026
600c67d2
88696c8c
40068d2d
3f3c4037
4f5c1040
433c0001
414c805e
23c3886c
46646026
08564196
00000804
bf961016
612c1364
32c34c09
0001341c
80378026
67d223c3
6c8c600c
10c3235c
60376006
10403f3c
00014f5c
805e433c
000e235c
886c414c
606623c3
41964664
08040856
bf961016
612c1364
34c38c09
0001341c
80378026
600c69d2
425c6c8c
435c001b
400610c6
3f3c4037
4f5c1040
433c0001
414c805e
23c3886c
46646026
08564196
00000804
bf96f016
71c350c3
625c7364
612c001b
31c32c09
0001341c
202623c3
60072037
800c1654
6d4c720c
366416c3
326430c3
20464006
331c2037
095400ff
0487333c
6d00502c
4eeb6c4c
60376006
10403f3c
00011f5c
805e133c
000e635c
001e235c
886c554c
17c305c3
60a623c3
41964664
08040f56
0136f016
50c3bf96
81c362c3
725c8364
612c001b
31c32c09
0001341c
40374026
1c546007
720c800c
17c36d4c
30c33664
20463264
331c2037
105400ff
0487333c
6c80302c
36c34c4c
02be133c
2c0b2aee
2717313c
40066a6f
3f3c4037
1f5c1040
133c0001
735c805e
554c000e
05c3886c
23c318c3
46646066
80764196
08040f56
0136f016
50c3bf96
81c372c3
625c8364
612c001b
31c32c09
0001341c
402666f2
43c34037
01f323c3
720c800c
16c36d4c
20c33664
323c2264
7fe50ff6
133c7f32
2037080c
10403f3c
00010f5c
805e033c
000e635c
2ff22017
0487323c
6d00502c
1ca96c8c
2ca905f2
003d1f5c
4ce90093
003d2f5c
8c6c754c
18c305c3
00402f3c
46646086
80764196
08040f56
bf96f016
71c350c3
625c7364
612c001b
31c32c09
0001341c
202623c3
60072037
800c1754
6d4c720c
366416c3
326430c3
20464006
331c2037
0a5400ff
0487333c
6d00502c
235c6c4c
60060233
3f3c6037
1f5c1040
133c0001
635c805e
235c000e
554c001e
05c3886c
23c317c3
466460a6
0f564196
00000804
0336f016
50c3be96
91c372c3
825c9364
612c001b
31c32c09
0001341c
40374026
28546007
d20c800c
18c3794c
30c33664
60773264
60376046
21c32057
00ff231c
20571954
0487313c
4c80302c
6d49682c
20372186
0e946047
275c684c
235c002b
78ac0236
2f5c05c3
12c30021
60063664
3f3c6037
1f5c1080
133c0001
835c805e
554c000e
05c3886c
23c319c3
46646066
c0764296
08040f56
bf963016
8c09612c
361c34c3
433c0001
80370014
00015f5c
00255f5c
8c69622c
002d4f5c
8c6c614c
00402f3c
46646046
0c564196
00000804
be961016
612c1364
32c34c09
0001341c
40374026
67d26077
6d4c600c
60776c69
60376006
00012f5c
00452f5c
00213f5c
004d3f5c
8c6c614c
00802f3c
46646046
08564296
00000804
bf961016
612c1364
34c38c09
0001341c
80378026
600c67d2
88696d4c
40068c6d
3f3c4037
4f5c1040
433c0001
414c805e
23c3886c
46646026
08564196
00000804
be961016
612c1364
32c34c09
0001341c
40374026
67d26077
6d0c600c
60776d09
60376006
00012f5c
00452f5c
00213f5c
004d3f5c
8c6c614c
00802f3c
46646046
08564296
00000804
bf961016
612c1364
34c38c09
0001341c
80378026
600c67d2
88696d0c
40068d0d
3f3c4037
4f5c1040
433c0001
414c805e
23c3886c
46646026
08564196
00000804
be961016
612c1364
32c34c09
0001341c
40374026
67d26077
6d8c600c
60776c89
60376006
00012f5c
00452f5c
00213f5c
004d3f5c
8c6c614c
00802f3c
46646046
08564296
00000804
bf961016
612c1364
34c38c09
0001341c
80378026
600c67d2
88696d8c
40068c8d
3f3c4037
4f5c1040
433c0001
414c805e
23c3886c
46646026
08564196
00000804
be967016
61c350c3
125c6364
612c001b
32c34c09
0001341c
40374026
18546007
8e0c600c
3664714c
326430c3
60466077
40576037
331c32c3
0a5400ff
05c3718c
00212f5c
366412c3
326430c3
3f3c6037
2f5c1080
233c0001
554c805e
05c3888c
23c316c3
46646026
0e564296
00000804
be967016
a809412c
361c35c3
533c0001
a0770014
00216f5c
00456f5c
623268a9
0014533c
6f5ca037
6f5c0001
614c004d
2f3c8c6c
60460080
42964664
08040e56
bd967016
61c350c3
012c6364
313c2009
80260014
600780b7
42c31d54
019e343c
67d240a9
627232c3
2f5c6077
00d30021
629232c3
2f5c6037
40ad0001
6e0c740c
6d6c546c
0110023c
36645009
326430c3
3f3c60b7
4f5c10c0
433c0041
554c805e
05c3886c
23c316c3
46646026
0e564396
00000804
be961016
612c1364
32c34c09
0001341c
40266037
67d24077
6c8c600c
60376ec8
60776006
00212f5c
00452f5c
00013f5c
004d3f5c
8c6c614c
00802f3c
46646046
08564296
00000804
bf963016
612c1364
34c38c09
0001341c
822c6fd2
600770a8
70880b74
08d46007
6c8c600c
aecda869
40374006
60260073
3f3c6037
4f5c1040
433c0001
414c805e
23c3886c
46646026
0c564196
00000804
be96f016
62c350c3
736471c3
001b125c
4c09612c
341c32c3
40260001
60074077
800c2054
6d4c720c
30c33664
40463264
331c4077
155400ff
0487333c
6d00502c
d8a96c4c
2f5cc037
235c0001
4226014d
40174077
402646f2
0155235c
60776017
10803f3c
00212f5c
805e233c
888c554c
17c305c3
602623c3
42964664
08040f56
0136f016
50c3be96
81c362c3
725c8364
612c001b
31c32c09
0001341c
40374026
60076077
800c2054
6d4c720c
366417c3
326430c3
20372046
40774006
00ff331c
333c1254
502c0487
4c8c6d00
602778a9
48e90694
40064077
00b34037
407748a9
60376006
10803f3c
00011f5c
805e133c
000e735c
00212f5c
005d2f5c
1f5c12c3
2f5c0065
554c006d
05c3886c
23c318c3
466460c6
80764296
08040f56
be963016
8006612c
00454f5c
45c3aca9
0001441c
5f5c8077
5f5c0021
6ca9004d
533c6132
a0370014
00013f5c
00553f5c
8c6c614c
00802f3c
46646066
0c564296
00000804
bf961016
612c1364
32c34c09
0001341c
802623c3
66d28037
6d6c600c
60064ccb
3f3c6037
4f5c1040
433c0001
235c805e
414c000e
23c3886c
46646066
08564196
00000804
bf961016
612c1364
34c38c09
0001341c
80378026
600c68d2
425c6d6c
8cce001b
40374006
10403f3c
00014f5c
805e433c
886c414c
602623c3
41964664
08040856
bf961016
612c1364
32c34c09
0001341c
80378026
66d223c3
6d0c600c
60064cab
3f3c6037
4f5c1040
433c0001
235c805e
414c000e
23c3886c
46646066
08564196
00000804
bf961016
612c1364
34c38c09
0001341c
80378026
600c68d2
425c6d0c
8cae001b
40374006
10403f3c
00014f5c
805e433c
886c414c
602623c3
41964664
08040856
c0967016
61c350c3
28696364
52bc4889
2f3c0943
60061000
805e323c
8c6c754c
16c305c3
60262fc3
40964664
08040e56
be96f016
52c360c3
736471c3
4c09612c
341c32c3
40260001
60074037
600c1a54
71ac8e0c
0030153c
30c33664
60773264
60376186
32c34057
00ff331c
70ec0a54
2f5c06c3
12c30021
36645529
60376006
10804f3c
00012f5c
805e243c
00900f3c
0030153c
094282bc
ac6c794c
17c306c3
60e624c3
42965664
08040f56
b7967016
61c350c3
612c6364
32c34c09
0001341c
40374026
600c69d2
6ccc6e0c
10401f3c
60063664
2f5c6037
2f5c0001
0f3c0025
1f3c0050
44061040
08cbb0bc
8c6c754c
16c305c3
00402f3c
46646426
0e564996
00000804
bf967016
61c350c3
612c6364
32c34c09
0001341c
40374026
10546007
6c8c600c
2f5c4e29
0f3c002d
133c0060
201c1270
b0bc00f0
600608cb
3f3c6037
2f5c1040
233c0001
554c805e
05c3886c
23c316c3
46647e46
0e564196
00000804
bf967016
61c350c3
612c6364
32c34c09
0001341c
40374026
600c6cd2
0f3c6c8c
133c0060
40660170
08cbb0bc
60376006
00012f5c
00252f5c
4c69762c
002d2f5c
8c6c754c
16c305c3
00402f3c
466460a6
0e564196
00000804
bf967016
61c350c3
612c6364
31c32c09
0001341c
20372026
600c6cd2
033c6c8c
123c0290
40660030
08cbb0bc
40374006
10403f3c
00011f5c
805e133c
886c554c
16c305c3
602623c3
41964664
08040e56
bf967016
61c350c3
612c6364
32c34c09
0001341c
40374026
600c6cd2
0f3c6c8c
133c0050
40660290
08cbb0bc
60376006
10403f3c
00012f5c
805e233c
886c554c
16c305c3
608623c3
41964664
08040e56
0f36f016
50c3b796
b1c302c3
752cb364
31c32c09
0001341c
40774026
600760b7
740c3954
cc8c4e10
0019905c
5889762c
403c6c49
20060040
207720b7
201423e4
08c30533
82bc14c3
07c30942
0060143c
b0bc4206
2ac308cb
05c3684c
27c318c3
60973664
202513c3
2f5c2037
40b70001
762c82c5
6c495889
061423e4
8f3c0133
7f3c11e0
409710e0
39e432c3
2006db14
2f5c2077
2f5c0021
3f5c0075
3f5c0041
754c007d
05c38c6c
2f3c1bc3
604600e0
49964664
0f56f076
00000804
0136f016
60c3be96
81c372c3
612c8364
32c34c09
0001341c
00770026
25546007
ac8c780c
564d4026
762d7c69
1270453c
101c04c3
9cbc00f0
04c308cb
0040173c
00f0201c
08cbb0bc
2160153c
00534006
32c44025
1dd205a2
6d207e06
2f5c6037
566d0001
60776006
10803f3c
00210f5c
805e033c
886c594c
18c306c3
602623c3
42964664
0f568076
00000804
c096f016
71c350c3
612c7364
32c34c09
0001341c
00106f3c
11546007
8c8c600c
3f5c6006
06c30005
02f0143c
b0bc5049
504908cb
40067900
01334c0d
3f5c6026
06c30005
00f8101c
08cb9cbc
8c6c754c
17c305c3
7f262fc3
40964664
08040f56
0f36f016
60c3bd96
b1c342c3
612cb364
31c32c09
0001341c
40374026
600723c3
a00c2b54
f48c1610
10609f3c
143c09c3
82bc0030
a75c0942
91290021
624686d2
80276037
01131494
686c28c3
19c306c3
80373664
7a2c0193
4c4915ec
0187123c
08cb9cbc
7c8d6006
20372006
3c892ac3
23c368a0
3f5c2364
3f5c0001
3f3c0035
235c0060
594c000e
06c3886c
23c31bc3
46646066
f0764396
08040f56
bf96f016
71c360c3
612c7364
31c32c09
0001341c
20372026
12546007
ac8c600c
0170453c
123c04c3
40660040
08cbb0bc
153c04c3
00bc2220
40060942
3f3c4037
1f5c1040
133c0001
594c805e
06c3886c
23c317c3
46646026
0f564196
00000804
efc34036
1f36f016
50c3bd96
b364b1c3
612ccfc3
31c32c09
0001341c
1e5c2026
13c3f6a7
54546007
c00cafc3
f88c1a10
2c49622c
0067313c
341c60c5
f3a40ffc
89299fc3
424688d2
f6a72e5c
80272006
02733e94
0030623c
65cc18c3
366416c3
32540007
682c28c3
202605c3
366426c3
f6a74e5c
05732026
7c898006
12946007
343c0473
243c0067
19c30187
79ec0580
82bc2980
243c0942
2e5c0010
4e5cf687
7c89f681
f6c73e5c
ec1443e4
682c28c3
2e5c05c3
12c3f6c1
366429c3
60063c89
f6a73e5c
20060093
f6a71e5c
2e3cfac3
3e5cfdc0
323cf6a1
762c805e
325c6c49
125c000e
754c001e
05c38c6c
60a61bc3
fcc34664
f8764396
ef3c0f56
0804024f
fe961016
226440c3
60373264
2c09612c
341c31c3
60070001
323c1754
60070014
614c1354
1f3c6e6c
5fe60040
40263664
1f5c400d
204d0001
714c402d
04c36c0c
40662057
02963664
08040856
fe967016
61c340c3
22646264
612c4037
31c32c09
0001341c
25546007
60aca00c
32c34c09
0020341c
1d546007
6e6c614c
00401f3c
36645fe6
600d60c6
00011f5c
363c204d
342c0487
6c2c6c80
0333135c
001e105c
602d6066
6c0c714c
205704c3
366440a6
0e560296
00000804
fe967016
61c340c3
22646264
612c4037
31c32c09
0001341c
25546007
60aca00c
32c34c29
0001341c
1d546007
6e6c614c
00401f3c
36645fe6
600d6126
00011f5c
363c204d
342c0487
6c2c6c80
0333135c
001e105c
602d6066
6c0c714c
205704c3
366440a6
0e560296
00000804
fe963016
126440c3
40372264
4c09612c
341c32c3
60070001
400c2954
0487313c
6c80282c
60acac2c
32c34c69
0008341c
1c546007
6e6c614c
00401f3c
36645fe6
200d2386
00012f5c
155c404d
105c0333
255c001e
205c0343
20a6002e
714c202d
04c36c0c
40e62057
02963664
08040c56
0736f016
50c3fd96
22641264
612c4077
32c34c09
0001341c
4e546007
813cc00c
782c0487
8d4c3884
2ca960ac
341c31c3
60070020
614c4154
1f3c6e6c
5fe60080
f14b3664
00b3945c
50c930a9
093412e4
3210141d
128da33c
0007af5c
00012f5c
200d25c6
00213f5c
782c604d
6c2c3884
0333635c
001e605c
61c330a9
363c30eb
305c128d
d0eb002e
628d323c
003e305c
105c312b
19c3004e
236429c3
023427e4
105c17c3
c166005e
754cc02d
05c36c0c
41a62097
03963664
0f56e076
00000804
ff967016
61c340c3
612c6264
31c32c09
0001341c
24546007
60aca00c
60076cc8
614c1f15
1fc36e6c
36645fe6
670620c3
163c600d
742c0487
6c2c6c80
0333035c
742c082e
6c4c6c80
0233135c
6086284e
714c682d
04c36c0c
40c62017
01963664
08040e56
fd967016
61c340c3
22646364
32644077
5f5c6037
60ac00e3
32c34c49
0008341c
1a546007
6e6c614c
00801f3c
36645fe6
400d4286
00212f5c
605c404d
2f5c001e
40ad0001
40c6a06e
714c402d
04c36c0c
41062097
03963664
08040e56
ff967016
61c340c3
22646264
0c09612c
341c30c3
60070001
30ac3254
0116323c
533c7fe5
0449f88c
341c30c3
62d20001
04e9a9f2
341c30c3
60070001
47272054
714c1e94
04c36e6c
5fe61fc3
a4d23664
400d4226
67260073
500c600d
0487363c
6c80282c
235c6c2c
402e0333
602d6046
6c0c714c
201704c3
36644086
0e560196
00000804
fe96f016
126460c3
40372264
4c09612c
341c32c3
60070001
400c2d54
0487313c
6c80282c
60acec2c
32c34c49
0002341c
20546007
614cbd49
1f3c6e6c
5fe60040
40c33664
600d6246
00011f5c
0065204d
82bc17c3
353c0942
33c40026
345c7f32
4106004f
794c502d
06c36c0c
41462057
02963664
08040f56
fe96f016
71c350c3
22647264
c00c4037
2c09612c
341c31c3
60070001
60ac2654
32c34ce9
0008341c
1f546007
6e6c614c
00401f3c
36645fe6
30c340c3
133c2786
273c015f
382c0487
03c34880
82bc282c
2f5c0942
510d0001
702d60e6
6c0c754c
205705c3
36644126
0f560296
00000804
fe96f016
61c370c3
612c6264
32c34c09
0001341c
2c546007
60aca00c
32c34ce9
0004341c
24546007
0487663c
6f00742c
60376c2c
6e6c614c
00401f3c
36645fe6
30c340c3
233c4766
03c3015f
82bc2017
742c0942
6c6c6f00
07a4235c
6146504f
7d4c702d
07c36c0c
41862057
02963664
08040f56
fe96f016
71c350c3
22647264
612c4037
32c34c09
0001341c
25546007
60acc00c
32c34cc9
0020341c
1d546007
6e6c614c
00401f3c
36645fe6
66c640c3
2f5c600d
404d0001
0487373c
6d00582c
2c2c0065
094282bc
702d60e6
6c0c754c
205705c3
36644126
0f560296
00000804
ff96f016
71c350c3
612c7264
31c32c09
0001341c
23546007
60acc00c
32c34cc9
0010341c
1b546007
6e6c614c
5fe61fc3
40c33664
26a630c3
015f133c
0487273c
4880382c
282c03c3
094282bc
502d40c6
6c0c754c
201705c3
36644106
0f560196
00000804
ff96f016
71c350c3
612c7264
31c32c09
0001341c
23546007
60acc00c
32c34cc9
0008341c
1b546007
6e6c614c
5fe61fc3
40c33664
268630c3
015f133c
0487273c
4880382c
282c03c3
094282bc
502d40c6
6c0c754c
201705c3
36644106
0f560196
00000804
0136f016
50c3ff96
71c382c3
612c7264
31c32c09
0001341c
24546007
60acc00c
32c34cc9
0004341c
1c546007
6e6c614c
5fe61fc3
40c33664
266630c3
015f133c
0487273c
4880382c
282c03c3
094282bc
41461051
754c502d
05c36c0c
41862017
01963664
0f568076
00000804
ff967016
126460c3
4c09612c
341c32c3
60070001
400c2a54
8cc960ac
341c34c3
60070002
313c2254
282c0487
ac2c6c80
6e6c614c
5fe61fc3
40c33664
464630c3
015f233c
15c303c3
094282bc
710d76e9
312d3709
514d5729
702d6126
6c0c794c
201706c3
36644166
0e560196
00000804
ff967016
126460c3
4c09612c
341c32c3
60070001
400c2454
8cc960ac
341c34c3
60070001
313c1c54
282c0487
ac2c6c80
6e6c614c
5fe61fc3
40c33664
462630c3
015f233c
15c303c3
094282bc
702d60c6
6c0c794c
201706c3
36644106
0e560196
00000804
ff967016
51c360c3
4c09612c
341c32c3
60070001
60ac2b54
32c34c89
0002341c
24546007
6e6c614c
5fe61fc3
40c33664
600d6446
404d4026
153c0065
82bc0010
74e90942
5509712d
7529516d
5549718d
752b51ad
540970ee
61e6520d
794c702d
06c36c0c
42262017
01963664
08040e56
ff96f016
71c350c3
612c7264
31c32c09
0001341c
23546007
60acc00c
32c34c49
0040341c
1b546007
6e6c614c
5fe61fc3
40c33664
22e630c3
015f133c
0487273c
4880382c
282c03c3
094282bc
502d40c6
6c0c754c
201705c3
36644106
0f560196
00000804
ff96f016
71c350c3
612c7264
31c32c09
0001341c
23546007
60acc00c
32c34c49
0020341c
1b546007
6e6c614c
5fe61fc3
40c33664
22c630c3
015f133c
0487273c
4880382c
282c03c3
094282bc
502d40c6
6c0c754c
201705c3
36644106
0f560196
00000804
ff967016
51c360c3
4c09612c
341c32c3
60070001
60ac2c54
32c34c09
0002341c
25546007
6e6c614c
5fe61fc3
40c33664
600d6046
404d4026
153c0065
82bc0010
74e90942
4006712d
750950ae
5529718d
754951ad
552b71cd
007e245c
702d61e6
6c0c794c
201706c3
36644226
0e560196
00000804
ff967016
126450c3
4c09612c
341c32c3
60070001
400c2b54
0487313c
6c80282c
60accc2c
32c34ce9
0010341c
1e546007
6e6c614c
5fe61fc3
40c33664
27a630c3
015f133c
16c303c3
094282bc
0080043c
0220163c
b0bc4106
41c608cb
754c502d
05c36c0c
42062017
01963664
08040e56
fe96f016
126450c3
40372264
4c09612c
341c32c3
60070001
400c2d54
0487313c
cc80282c
60acf82c
60076c48
614c2315
1f3c6e6c
5fe60040
40c33664
230630c3
015f133c
17c303c3
094282bc
043c786c
133c0080
420600e0
08cbb0bc
00012f5c
62e6530d
754c702d
05c36c0c
43262057
02963664
08040f56
fe967016
126450c3
40372264
4c09612c
341c32c3
60070001
400c2c54
0487313c
6c80282c
60accc2c
32c34c29
0004341c
1f546007
6e6c614c
00401f3c
36645fe6
616640c3
1f5c600d
204d0001
0333265c
001e205c
163c00a5
410601a0
08cbb0bc
702d6166
6c0c754c
205705c3
366441a6
0e560296
00000804
fe967016
126450c3
40372264
4c09612c
341c32c3
60070001
400c3954
0487313c
6c80282c
60accc2c
32c34c09
0040341c
24546007
6e6c614c
00401f3c
36645fe6
60e640c3
1f5c600d
204d0001
16c30065
094282bc
0090043c
5a89388c
08cbb0bc
71005a89
2d2d2006
502d5fe6
6c0c754c
205705c3
0101201c
388c3664
758c27d2
05c36c2c
60063664
0296788f
08040e56
fc967016
31c350c3
60b73264
40772264
4c09612c
341c32c3
60070001
200c3f54
343c8097
842c0487
c82c4e00
8c0960ac
341c34c3
60370008
23546007
6e6c614c
00c01f3c
36645fe6
30c340c3
233c4086
03c3015f
82bc16c3
043c0942
163c0080
406600b0
08cbb0bc
00213f5c
4146716d
754c502d
05c36c0c
418620d7
01d33664
6beb484c
6bee6072
6d0c660c
00414f5c
4f5c14c3
24c30001
04963664
08040e56
ff967016
51c360c3
4c09612c
341c32c3
60070001
60ac4354
32c34ca9
0040341c
3c546007
6e6c614c
5fe61fc3
40c33664
600d65e6
404d4026
153c0065
82bc0010
74e90942
5509712d
7529516d
5549718d
752b51ad
540970ee
346c520d
231c5609
033500ef
00f0201c
0110043c
08cbb0bc
301c3609
4ca000f0
07f44007
0110313c
12c31180
08cb9cbc
502d5fe6
6c0c794c
201706c3
0101201c
01963664
08040e56
0136f016
80c3fc96
52c331c3
60b73264
2c4960ac
341c31c3
60070010
614c3754
1f3c6e6c
5fe600c0
70c33664
400d42a6
00413f5c
403c604d
65c30030
0253a006
16c304c3
b0bc40c6
043c08cb
22060060
08cb9cbc
0010253c
5f5c4077
82c50021
6097c0c5
51e413c3
333cec14
233c0167
123c0030
2037ffe0
00013f5c
18c37c2d
6c0c654c
20d708c3
04963664
0f568076
00000804
fe967016
126460c3
40372264
4c09612c
341c32c3
60070001
400c3454
0487313c
6c80282c
60acac2c
32c34c29
0010341c
27546007
6e6c614c
00401f3c
36645fe6
61a640c3
1f5c600d
204d0001
0333255c
001e205c
60ad6006
20cd3509
210600e5
08cb9cbc
245c57cc
7fe6007f
009f345c
302d22a6
6c0c794c
205706c3
366442e6
0e560296
00000804
fd967016
126460c3
22642077
60373264
323c200c
442c0487
ac2c6d00
4c8960ac
341c32c3
60070004
1f3c3854
5fe60080
094488bc
646640c3
2f5c600d
404d0021
0333355c
001e305c
00012f5c
355c40ad
60cd0191
45f24017
153c00e5
011301a0
23c36017
08944027
153c00e5
41060220
08cbb0bc
00e50173
23c36017
02a0153c
f6544047
9cbc2106
61a608cb
06c3702d
41e62097
09466abc
0e560396
00000804
0336f016
50c3ff96
226421c3
2c09612c
341c31c3
60070001
c00c3454
0487323c
582c93c3
39c39284
60acec2c
31c32c69
0004341c
25546007
6e6c614c
5fe61fc3
40c33664
400d4366
0333375c
175c602e
208d01c1
784c1890
444c19c3
125c0e69
275c0203
e0bc01c1
28c30986
1106025c
702d6066
6c0c754c
201705c3
366440a6
c0760196
08040f56
ff961016
326431c3
000c6037
6aa9408c
41c32017
125434e4
f5242e24
00013f5c
80176aad
402724c3
412c0594
8fcc60ec
313c884f
62d24004
0196f324
08040856
1f36f016
41c3fe96
612c4364
32c34c09
0001341c
53546007
ae246010
622cf524
0001a35c
094b343c
0287933c
098b343c
0347833c
60776006
743c03c3
643c0104
06b30804
682c2bc3
442c2c00
602768e9
68c92694
23546007
0333325c
079434e4
4004353c
2e546007
0593f324
64ececd2
6d893984
13946027
4004353c
22546007
0413f324
64ccccd2
6d2228c3
07946027
4004353c
16546007
0293f324
32c34057
60376025
00012f5c
09054077
c3c36057
c914cae4
4004353c
f32462d2
00ff301c
2f5c6077
02c30021
f8760296
08040f56
ff967016
d48ca00c
6dcc760c
00073664
8e241654
5889f524
0187323c
2d0055ec
b0bc4306
788908cb
5fe523c3
3f5c4037
788d0001
4004343c
f32462d2
0e560196
00000804
3f36f016
b0c3ff96
326431c3
042c200c
0487333c
48304180
c86ce84c
64aca890
313c2c29
81800487
30301050
9090b06c
652c1bc3
23722ca9
1f5c2037
2cad0001
1ac36026
2006652d
1ac33f6d
01c5315c
0380023c
0380143c
e6bc4186
b01c08cb
71f10000
71d17211
4beb28c3
39c35fee
01a1135c
135c3ac3
28c301a5
5ecf4acc
6fcb38c3
18c37fce
3eef26ec
490928c3
38c35d0d
7d2d6d29
670c18c3
7f0f6a92
590d5509
0203315c
0206375c
3dcd25c9
49e928c3
38c35ded
7e0d6e09
215c19c3
1ac30333
0336215c
6e8939c3
19c3668d
0191215c
215c1ac3
39c30195
66ed6ee9
470919c3
470d1ac3
6f2939c3
063c672d
153c00e0
420600e0
08cbb0bc
01e0063c
01e0153c
b0bc4206
063c08cb
153c02e0
420602e0
08cbb0bc
03e0063c
03e0153c
b0bc4206
063c08cb
153c0b60
46060b60
08cbb0bc
05e0063c
05e0153c
b0bc4206
063c08cb
153c06e0
420606e0
08cbb0bc
07e0063c
07e0153c
b0bc4206
063c08cb
153c09e0
430609e0
08cbb0bc
08e0063c
08e0153c
b0bc4206
0a3c08cb
193c01a0
410601a0
08cbb0bc
02200a3c
0220193c
b0bc4106
19c308cb
1ac3448c
39c3448f
34496c91
255c384d
265c07a4
74c907a7
34e978cd
552938ed
38c3592d
7f8e6f8b
394d3549
596d5569
798d7589
215c19c3
1ac303a3
03a6215c
6fe938c3
18c37fed
0233115c
0236175c
4ae928c3
3cc35eed
3dc32c69
2cc32c6d
4c8d4889
2d093cc3
2d0d3dc3
586d5469
788d7489
38ad34a9
04e0063c
04e0153c
b0bc4206
28c308cb
5d8d4989
fc760196
08040f56
0136f016
60c3ff96
72c381c3
b08c800c
6dcc720c
07d23664
17c300c5
b0bc4206
03f308cb
7a2c5489
32e46c49
323c1a35
51ec0187
18c30d00
094282bc
313c3489
51ec0187
033c6d00
17c30060
b0bc4206
748908cb
202513c3
2f5c2037
548d0001
80760196
08040f56
fe96f016
71c340c3
2c09612c
341c31c3
60070001
c00c3354
f524ae24
03f34006
313c2057
582c0487
2c2c6d00
600764c9
64e91054
0d946027
88bc07c3
30c30942
67f23264
4004353c
1b546007
0333f324
13c36057
20372025
00012f5c
722c4077
20576c09
32e421c3
353cdcb4
66d24004
101cf324
207700ff
301c0093
607700ff
00211f5c
029601c3
08040f56
51c37016
63c342c3
60476549
116f1294
345c6069
606901e5
400673ee
0185245c
01cd245c
24bc02c3
063c094a
023322a0
6469316f
01e5345c
73ee6469
245c4026
245c0185
02c301cd
094a24bc
05e0053c
01e1145c
01f1245c
097bfebc
345c6006
345c012d
345c0135
0e56018d
00000804
fe967016
226441c3
606c4077
716f200c
245c4c69
6c6901e5
73ee6037
645cc006
a026012d
645cb20d
545c0135
545c0185
648c018d
22a0033c
3f5c12c3
23c30001
097bfebc
3f5c05c3
13c30021
d6bc24c3
06c3094a
01c9145c
094ba4bc
0e560296
00000804
ff96f016
226441c3
616c4037
323c4c69
402c0487
cc2c6d00
7869c56f
01e5315c
67ee7869
715ce026
715c012d
a0060135
0185515c
01cd515c
018d515c
24bc05c3
063c094a
145c05e0
245c01e1
febc01f1
07c3097b
00012f5c
24c312c3
094ad6bc
145c05c3
a4bc01c9
0196094b
08040f56
ff967016
226441c3
608c4037
656f62e5
615cc006
400601e5
215c47ee
a026012d
615ca60d
515c0135
515c0185
608c018d
2220033c
febc16c3
05c3097b
00013f5c
24c313c3
094ad6bc
145c06c3
a4bc01c9
0196094b
08040e56
ff96f016
41c370c3
40372264
63a5608c
a006656f
01e5515c
67ee6006
615cc026
615c012d
315c0135
515c0185
515c01cd
6006018d
05c3646f
094a24bc
033c7c8c
145c2220
245c01e1
febc01f1
05c3097b
00013f5c
24c313c3
094ad6bc
145c06c3
a4bc01c9
0196094b
08040f56
50c33016
405c8006
405c01cd
405c0135
405c012d
405c0185
04c3018d
094a24bc
155c04c3
a4bc01c9
0c56094b
00000804
fb961016
105c2026
2f3c01dd
101c0140
123c0c03
2006fe6e
00951f5c
3f3c200c
60370130
3f5c6026
3f3c0025
60b700c0
101c840c
60660c03
00d74664
3f5c05f2
62d20099
059603c3
08040856
f896f016
01a36f5c
405c8026
4f3c01dd
701c0200
743c0c33
e0e6f76e
00857f5c
001e145c
009d2f5c
d08e706e
3f3c400c
603701f0
3f5c6026
3f3c0025
60b70180
101ca80c
24c30c33
56646146
05f20197
00f93f5c
03c362d2
0f560896
00000804
0136f016
61c3f896
83c372c3
205c4026
2f3c01dd
301c0200
323c1005
6006feee
00fd3f5c
5f3c200c
a03700e0
3f5c6146
3f3c0025
60b70180
101c840c
60661005
01974664
12940007
00713f5c
03c363d2
255c01b3
580e000b
00893f5c
544b7c0e
4c0e38c3
6397546b
08964c0e
0f568076
00000804
f6961016
20262177
01dd105c
02802f3c
0c24401c
f96e423c
1f5c2066
4f5c00e5
4f5c00a1
215700ed
420b413c
4f5c8137
4f5c0081
215700f5
440b413c
4f5c80f7
4f5c0061
200c00fd
02703f3c
60266037
00253f5c
02003f3c
840c60b7
0c24101c
466460c6
05f20217
01393f5c
03c362d2
08560a96
00000804
f7963016
402652c3
01dd205c
02402f3c
1405401c
f5ee423c
4f5c8046
125c008d
200c001e
01c03f3c
60866037
00253f5c
02003f3c
840c60b7
1405101c
466460a6
69f26217
00e13f5c
68f203c3
00f94f5c
0073940d
540d4006
09960217
08040c56
f9967016
402662c3
01dd205c
01c02f3c
0c7b401c
fbee423c
4f5c8046
125c00ad
200c001e
00e05f3c
60a6a037
00253f5c
01803f3c
840c60b7
0c7b101c
466460a6
09f20197
00713f5c
03c363d2
455c0093
980e001b
0e560796
00000804
f9963016
405c8026
4f3c01dd
501c01c0
543c0c7c
a086f86e
00755f5c
001e145c
002e245c
3f3c400c
60370130
3f5c6066
3f3c0025
60b70180
101ca80c
24c30c7c
566460e6
05f20197
00993f5c
03c362d2
0c560796
00000804
f8961016
402640f7
01dd205c
02002f3c
0406401c
f96e423c
4f5c8066
125c00a5
1f5c001e
1f5c0061
200c00bd
01f03f3c
60266037
00253f5c
01803f3c
840c60b7
0406101c
466460c6
05f20197
00f93f5c
03c362d2
08560896
00000804
f9963016
402652c3
01dd205c
01c02f3c
1403401c
f9ee423c
4f5c8046
125c008d
200c001e
01403f3c
60866037
00253f5c
01803f3c
840c60b7
1403101c
466460a6
69f26197
00a13f5c
68f203c3
00b94f5c
0073940d
540d4006
07960197
08040c56
f9963016
405c8026
4f3c01dd
501c01c0
543cfc06
a046f9ee
008d5f5c
00951f5c
009d2f5c
3f3c400c
603701b0
3f5c6026
3f3c0025
60b70140
101ca80c
24c3fc06
566460a6
05f20157
00d93f5c
03c362d2
0c560796
00000804
f8967016
602650c3
01dd305c
02004f3c
0c01301c
f6ee343c
3f5c6106
0f3c007d
41060100
08cbb0bc
3f3c540c
603701f0
3f5c6026
3f3c0025
60b70180
05c3c80c
0c01101c
616624c3
01976664
3f5c05f2
62d200f9
089603c3
08040e56
f8963016
202651c3
01dd105c
02002f3c
1009101c
feee123c
1f5c2006
200c00fd
00e03f3c
61466037
00253f5c
01803f3c
840c60b7
1009101c
46646066
6bf26197
00713f5c
68f203c3
1f3c05c3
40c600f0
08cbb0bc
08960197
08040c56
0136f016
60c3e396
82c371c3
03e05f3c
200605c3
bebc4646
4f3c0891
04c300c0
46462006
0891bebc
47374006
0c6c301c
2f5c740e
60260205
01dd365c
8037580c
3f5c6066
3f3c0025
60b70700
06c3880c
0c6c101c
606625c3
07174664
3f5c0df2
63d20061
011303c3
00692f5c
2f5c5c0d
38c30071
1d964c0d
0f568076
00000804
e1967016
126460c3
22642137
5f3c40f7
05c30460
46462006
0891bebc
01404f3c
200604c3
bebc4646
60060891
301c67b7
740e0c6d
3f5c6046
3f5c0245
3f5c0081
3f5c024d
3f5c0061
60260255
01dd365c
8037580c
00253f5c
07803f3c
880c60b7
101c06c3
25c30c6d
466460a6
05f20797
00a13f5c
03c362d2
0e561f96
00000804
0336f016
60c3e396
92c381c3
03e05f3c
200605c3
bebc4646
7f3c0891
07c300c0
46462006
0891bebc
47374006
2002301c
2f5c740e
60260205
01dd365c
e037580c
3f5c6086
3f3c0025
60b70700
06c3880c
2002101c
606625c3
07174664
3f5c0ef2
63d20061
013303c3
000b375c
680e28c3
00793f5c
680d29c3
c0761d96
08040f56
e396f016
71c350c3
03e06f3c
200606c3
bebc4646
4f3c0891
04c300c0
46462006
0891bebc
67376006
2007301c
6006780e
02053f5c
355c6026
540c01dd
60468037
00253f5c
07003f3c
880c60b7
101c05c3
26c32007
46646066
09f20717
00613f5c
03c363d2
3f5c0093
7c0d0069
0f561d96
00000804
e2967016
20f750c3
04206f3c
200606c3
bebc4646
4f3c0891
04c30100
46462006
0891bebc
67776006
200a301c
6026780e
02253f5c
00613f5c
022d3f5c
355c6026
540c01dd
3f5c8037
3f3c0025
60b70740
05c3880c
200a101c
608626c3
07574664
3f5c05f2
62d20081
1e9603c3
08040e56
e396f016
41c360c3
03e05f3c
200605c3
bebc4646
7f3c0891
07c300c0
46462006
0891bebc
67376006
200b301c
60e6740e
02053f5c
3f5c7009
702b020d
704b744e
70c9746e
02353f5c
3f5c7029
6026023d
01dd365c
e037580c
00253f5c
07003f3c
880c60b7
101c06c3
25c3200b
46646146
05f20717
00613f5c
03c362d2
0f561d96
00000804
e1967016
213760c3
5f3c40f7
05c30460
46462006
0891bebc
01404f3c
200604c3
bebc4646
60060891
301c67b7
740e200c
3f5c6046
3f5c0245
3f5c0081
3f5c024d
3f5c0061
60260255
01dd365c
8037580c
00253f5c
07803f3c
880c60b7
101c06c3
25c3200c
466460a6
05f20797
00a13f5c
03c362d2
0e561f96
00000804
e3967016
6f3c50c3
06c303e0
46462006
0891bebc
00c04f3c
200604c3
bebc4646
60060891
301c6737
780e200e
3f5c6006
60260205
01dd355c
8037540c
00253f5c
07003f3c
880c60b7
101c05c3
26c3200e
46646066
05f20717
00613f5c
03c362d2
0e561d96
00000804
e396f016
71c350c3
03e06f3c
200606c3
bebc4646
4f3c0891
04c300c0
46462006
0891bebc
67376006
200f301c
6006780e
02053f5c
355c6026
540c01dd
60468037
00253f5c
07003f3c
880c60b7
101c05c3
26c3200f
46646066
09f20717
00613f5c
03c363d2
3f5c0093
7c0d0069
0f561d96
00000804
e3967016
6f3c50c3
06c303e0
46462006
0891bebc
00c04f3c
200604c3
bebc4646
60060891
301c6737
780e2010
3f5c6006
60260205
01dd355c
8037540c
00253f5c
07003f3c
880c60b7
101c05c3
26c32010
46646066
05f20717
00613f5c
03c362d2
0e561d96
00000804
ef96f016
52c360c3
736471c3
00e04f3c
200604c3
bebc4646
60060891
101c6437
300e2013
3f5c61c6
745c0085
740b001e
002e345c
345c742b
744b003e
004e345c
345c746b
748b005e
006e345c
345c74ab
6026007e
01dd365c
6006580c
3f5c6037
3f3c0025
60b70400
06c3a80c
622624c3
04175664
0f561196
00000804
e396f016
71c360c3
4f3c7364
04c303e0
46462006
0891bebc
00c05f3c
200605c3
bebc4646
60060891
301c6737
700e201b
3f5c6046
745c0205
6026001e
01dd365c
a037580c
3f5c6066
3f3c0025
60b70700
06c3a80c
201b101c
60a624c3
07175664
3f5c05f2
62d20061
1d9603c3
08040f56
e2967016
126460c3
5f3c20f7
05c30420
46462006
0891bebc
01004f3c
200604c3
bebc4646
60060891
301c6777
740e201d
3f5c6026
3f5c0225
3f5c0061
6026022d
01dd365c
8037580c
00253f5c
07403f3c
880c60b7
101c06c3
25c3201d
46646086
05f20757
00813f5c
03c362d2
0e561e96
00000804
e0967016
126460c3
22642177
32644137
5f3c60f7
05c304a0
46462006
0891bebc
01804f3c
200604c3
bebc4646
60060891
301c67f7
740e201e
3f5c6066
3f5c0265
3f5c00a1
3f5c026d
3f5c0061
3f5c0275
3f5c0081
6026027d
01dd365c
8037580c
00253f5c
07c03f3c
880c60b7
101c06c3
25c3201e
466460c6
05f207d7
00c13f5c
03c362d2
0e562096
00000804
0136f016
50c3e396
6f3c81c3
06c303e0
46462006
0891bebc
00c07f3c
200607c3
bebc4646
40060891
301c4737
780e201f
02052f5c
355c6026
540c01dd
6066e037
00253f5c
07003f3c
880c60b7
101c05c3
26c3201f
46646066
0af20717
00613f5c
03c363d2
375c00b3
28c3000b
1d96680e
0f568076
00000804
0336f016
70c3e396
91c352c3
4f3c9364
c64603e0
200604c3
bebc26c3
8f3c0891
08c300c0
26c32006
0891bebc
67376006
2020101c
61c6300e
02053f5c
001e945c
345c740b
742b002e
003e345c
345c744b
746b004e
005e345c
345c748b
74ab006e
007e345c
375c6026
5c0c01dd
00078f5c
3f5c6066
3f3c0025
60b70700
07c3a80c
622624c3
07175664
c0761d96
08040f56
0136f016
60c3e296
836481c3
40f72264
04205f3c
05c38646
24c32006
0891bebc
01007f3c
200607c3
bebc24c3
40060891
101c4777
340e2021
3f5c6066
855c0225
2f5c001e
2f5c0061
4026023d
01dd265c
e037580c
00253f5c
07403f3c
880c60b7
25c306c3
466460c6
1e960757
0f568076
00000804
0336f016
60c3e396
736471c3
836482c3
936493c3
03e04f3c
200604c3
bebc4646
5f3c0891
05c300c0
46462006
0891bebc
67376006
2022101c
40c6300e
02052f5c
001e745c
002e845c
003e945c
365c6026
580c01dd
2066a037
00251f5c
07003f3c
a80c60b7
101c06c3
24c32022
56646126
05f20717
00613f5c
03c362d2
c0761d96
08040f56
0336f016
60c3e396
92c381c3
03e05f3c
200605c3
bebc4646
7f3c0891
07c300c0
46462006
0891bebc
47374006
2023301c
2f5c740e
60260205
01dd365c
e037580c
3f5c60a6
3f3c0025
60b70700
06c3880c
2023101c
606625c3
07174664
3f5c0ef2
63d20061
013303c3
000b375c
680e28c3
001b375c
680e29c3
c0761d96
08040f56
0136f016
60c3e396
736471c3
836482c3
03e04f3c
200604c3
bebc4646
5f3c0891
05c300c0
46462006
0891bebc
67376006
2024301c
6086700e
02053f5c
001e745c
002e845c
365c6026
580c01dd
3f5ca037
3f3c0025
60b70700
06c3a80c
2024101c
60e624c3
07175664
3f5c05f2
62d20061
1d9603c3
0f568076
00000804
e3967016
6f3c50c3
06c303e0
46462006
0891bebc
00c04f3c
200604c3
bebc4646
60060891
301c6737
780e2025
3f5c6006
60260205
01dd355c
8037540c
00253f5c
07003f3c
880c60b7
101c05c3
26c32025
46646066
05f20717
00613f5c
03c362d2
0e561d96
00000804
de96f016
71c350c3
00c06f3c
200606c3
bebc48c6
4f3c0891
04c30520
46462006
0891bebc
68776006
2026301c
6806780e
00753f5c
00f00f3c
480617c3
08cbb0bc
355c6026
540c01dd
3f5c8037
3f3c0025
60b70840
05c3880c
2026101c
686626c3
08574664
3f5c05f2
62d20291
229603c3
08040f56
e396f016
71c350c3
03e06f3c
200606c3
bebc4646
4f3c0891
04c300c0
46462006
0891bebc
67376006
201c301c
6006780e
02053f5c
355c6026
540c01dd
61268037
00253f5c
07003f3c
880c60b7
101c05c3
26c3201c
46646066
0cf20717
00613f5c
68f203c3
1f3c07c3
410600d0
08cbb0bc
1d960717
08040f56
0136f016
60c3e396
71c382c3
5f3c7364
05c303e0
46462006
0891bebc
00c04f3c
200604c3
bebc4646
60060891
301c6737
740e201a
3f5c6246
755c0205
0f3c001e
18c30430
b0bc4206
602608cb
01dd365c
8037580c
3f5c6066
3f3c0025
60b70700
06c3880c
201a101c
62a625c3
07174664
3f5c05f2
62d20061
1d9603c3
0f568076
00000804
0336f016
60c3e396
71c382c3
93c37364
5f3c9364
05c303e0
46462006
0891bebc
00c04f3c
200604c3
bebc4646
60060891
201c6737
540e2019
3f5c6386
755c0205
0f3c001e
18c30430
b0bc4106
955c08cb
0f3c006e
291704d0
b0bc4206
402608cb
01dd265c
8037580c
3f5c6026
3f3c0025
60b70700
06c3880c
2019101c
63e625c3
07174664
3f5c05f2
62d20061
1d9603c3
0f56c076
00000804
e396f016
71c350c3
03e06f3c
200606c3
bebc4646
4f3c0891
04c300c0
46462006
0891bebc
67376006
2018301c
6006780e
02053f5c
355c6026
540c01dd
61268037
00253f5c
07003f3c
880c60b7
101c05c3
26c32018
46646066
0cf20717
00613f5c
68f203c3
1f3c07c3
410600d0
08cbb0bc
1d960717
08040f56
0336f016
60c3e396
82c371c3
5f3c93c3
05c303e0
46462006
0891bebc
00c04f3c
200604c3
bebc4646
60060891
301c6737
740e2017
3f5c6406
0f3c0205
17c30410
b0bc4206
0f3c08cb
18c30510
b0bc4206
602608cb
01dd365c
8037580c
3f5c6226
3f3c0025
60b70700
06c3880c
2017101c
646625c3
07174664
3f5c0cf2
03c30061
09c368f2
00d01f3c
b0bc4206
071708cb
c0761d96
08040f56
e2967016
1f5c50c3
6f3c0076
06c30420
46462006
0891bebc
01004f3c
200604c3
bebc4646
60060891
301c6777
780e2016
3f5c6046
0f3c0225
1f3c0450
404600e0
08cbb0bc
355c6026
540c01dd
3f5c8037
3f3c0025
60b70740
05c3880c
2016101c
60a626c3
07574664
3f5c05f2
62d20081
1e9603c3
08040e56
0136f016
60c3e296
00761f5c
5f3c82c3
05c30420
46462006
0891bebc
01007f3c
200607c3
bebc4646
20060891
301c2777
740e2015
1f5c2046
0f3c0225
1f3c0450
404600e0
08cbb0bc
365c6026
580c01dd
2106e037
00251f5c
07403f3c
880c60b7
101c06c3
25c32015
466460a6
00070757
3f5c1594
03c30081
10946007
00732f5c
000b375c
099423e4
67d238c3
1f3c08c3
40a60130
08cbb0bc
1e960757
0f568076
00000804
e396f016
71c350c3
03e06f3c
200606c3
bebc4646
4f3c0891
04c300c0
46462006
0891bebc
67376006
2014301c
60a6780e
02053f5c
04100f3c
40a617c3
08cbb0bc
355c6026
540c01dd
3f5c8037
3f3c0025
60b70700
05c3880c
2014101c
610626c3
07174664
3f5c05f2
62d20061
1d9603c3
08040f56
e296f016
72c360c3
20f71264
04205f3c
200605c3
bebc4646
4f3c0891
04c30100
46462006
0891bebc
67776006
2012301c
60e6740e
02253f5c
00613f5c
022d3f5c
04600f3c
410617c3
08cbb0bc
365c6026
580c01dd
3f5c8037
3f3c0025
60b70740
06c3880c
2012101c
614625c3
07574664
3f5c05f2
62d20081
1e9603c3
08040f56
e296f016
72c360c3
20f71264
04205f3c
200605c3
bebc4646
4f3c0891
04c30100
46462006
0891bebc
67776006
2011301c
60e6740e
02253f5c
00613f5c
022d3f5c
04600f3c
410617c3
08cbb0bc
365c6026
580c01dd
3f5c8037
3f3c0025
60b70740
06c3880c
2011101c
614625c3
07574664
3f5c05f2
62d20081
1e9603c3
08040f56
e396f016
41c360c3
03e05f3c
200605c3
bebc4646
7f3c0891
07c300c0
46462006
0891bebc
47374006
200d301c
4326740e
02052f5c
355c70ab
50cb001e
002e255c
3f5c70e9
34c3022d
009f233c
02352f5c
04700f3c
40c613c3
08cbb0bc
3f5c7109
50eb026d
710b550e
512b752e
714b554e
516b756e
718b558e
402675ae
01dd265c
e037580c
3f5c6026
3f3c0025
60b70700
06c3880c
200d101c
638625c3
07174664
3f5c05f2
62d20061
1d9603c3
08040f56
e396f016
41c360c3
03e05f3c
200605c3
bebc4646
7f3c0891
07c300c0
46462006
0891bebc
67376006
2006301c
61e6740e
02053f5c
355c70ab
70cb001e
002e355c
3f5c7009
71c9022d
02353f5c
3f5c7049
0f3c023d
143c0480
40c60030
08cbb0bc
3f5c71e9
70290275
027d3f5c
365c6026
580c01dd
3f5ce037
3f3c0025
60b70700
06c3880c
2006101c
624625c3
07174664
3f5c05f2
62d20061
1d9603c3
08040f56
e396f016
71c350c3
03e06f3c
200606c3
bebc4646
4f3c0891
04c300c0
46462006
0891bebc
67376006
2005301c
60c6780e
02053f5c
04100f3c
410617c3
08cbb0bc
355c6026
540c01dd
3f5c8037
3f3c0025
60b70700
05c3880c
2005101c
612626c3
07174664
3f5c05f2
62d20061
1d9603c3
08040f56
e396f016
71c350c3
03e06f3c
200606c3
bebc4646
4f3c0891
04c300c0
46462006
0891bebc
67376006
2003301c
6006780e
02053f5c
355c6026
540c01dd
61268037
00253f5c
07003f3c
880c60b7
101c05c3
26c32003
46646066
0cf20717
00613f5c
68f203c3
1f3c07c3
410600d0
08cbb0bc
1d960717
08040f56
e396f016
71c350c3
03e06f3c
200606c3
bebc4646
4f3c0891
04c300c0
46462006
0891bebc
67376006
2001301c
6106780e
02053f5c
04100f3c
410617c3
08cbb0bc
355c6026
540c01dd
3f5c8037
3f3c0025
60b70700
05c3880c
2001101c
616626c3
07174664
3f5c05f2
62d20061
1d9603c3
08040f56
e196f016
71c360c3
000752c3
20075054
40074e54
40064c54
4f3c47b7
04c30460
464612c3
0891bebc
2009301c
4406700e
02452f5c
25c3a0f7
03f443e7
60f763e6
00612f5c
3f5c4137
3f5c0081
4f3c024d
04c30140
46462006
0891bebc
04605f3c
04a00f3c
411717c3
08cbb0bc
32c34117
15806085
2d2063e6
08cb9cbc
365c6026
580c01dd
3f5c8037
3f3c0025
60b70780
06c3880c
2009101c
646625c3
07974664
3f5c08f2
65d200a1
007303c3
0101001c
0f561f96
00000804
e196f016
71c360c3
000752c3
20075054
40074e54
40064c54
4f3c47b7
04c30460
464612c3
0891bebc
2008301c
4406700e
02452f5c
25c3a0f7
03f443e7
60f763e6
00612f5c
3f5c4137
3f5c0081
4f3c024d
04c30140
46462006
0891bebc
04605f3c
04a00f3c
411717c3
08cbb0bc
32c34117
15806085
2d2063e6
08cb9cbc
365c6026
580c01dd
3f5c8037
3f3c0025
60b70780
06c3880c
2008101c
646625c3
07974664
3f5c08f2
65d200a1
007303c3
0101001c
0f561f96
00000804
f8967016
02d242c3
001c24f2
06b30101
205c66c9
62c301d1
c077c025
00212f5c
6f5c40b7
605c0041
698001d5
2f5c6037
46cd0001
02003f3c
4d72458b
f66e233c
cc2ec206
4c4e4186
cc6ec0a6
2f5c4246
6f5c00a5
6f5c0001
410600ad
d00b4cae
502bccce
d04b4cee
506bcd0e
400c4d2e
13c3882c
46644286
0e560896
00000804
fc963016
536452c3
24f202d2
0101001c
3f3c0373
458b0100
233c4d72
4146f96e
40c64c2e
40a64c4e
42664c6e
00552f5c
2f5c4669
4046005d
acce4cae
882c400c
41c613c3
04964664
08040c56
fb961016
00e14f5c
4f3c8037
258b0140
143c2d72
2126f9ee
20a6302e
2086304e
2026306e
007d1f5c
00852f5c
3f5c70ae
3f5c0001
600c009d
14c36c2c
366441a6
08560596
00000804
fd967016
60ec51c3
04c3135c
236442c3
336431c3
023523e4
3f3c41c3
558b00c0
233c4d72
40e6faee
c0664c2e
4086cc4e
c0464c6e
004d6f5c
004e435c
882c400c
416613c3
03964664
08040e56
fd967016
60ec51c3
04c3135c
236442c3
336431c3
023523e4
3f3c41c3
558b00c0
233c4d72
40e6faee
c0664c2e
4086cc4e
6f5c4c6e
435c004d
400c004e
13c3882c
46644166
0e560396
00000804
fc961016
01004f3c
2d72258b
f9ee143c
302e2126
304e20a6
306e2086
005d1f5c
004e245c
005e345c
6c2c600c
41a614c3
04963664
08040856
50c3f016
62c341c3
73c36364
00077364
00ec2e54
04a4305c
29546007
27542007
6cac742c
3fe60c85
00073664
74ec2294
04a4335c
4d72518b
41264c0e
40a64c2e
40864c4e
40e64c6e
635c4d0d
735c004e
540c005e
05c3882c
41a613c3
742c4664
6cec54ec
0640023c
00733664
0101001c
08040f56
f8967016
c31750c3
43c32364
02d24364
001c24f2
06530101
02000f3c
6d72658b
f0ee303c
606e6086
3f5c6106
205c004d
405c004e
780c005e
06946047
305c784b
81e6006e
80060173
08946207
6c8c746c
00e00f3c
366416c3
14c383a6
2f3c1364
313c0010
682effc0
ff80313c
740c684e
05c36c2c
24c312c3
08963664
08040e56
fd961016
00c03f3c
2d72258b
faee133c
2c2e20e6
2c4e2066
2c6e2086
1f5c2146
235c004d
400c004e
13c3882c
46644166
08560396
00000804
fc961016
01004f3c
2d72258b
f9ee143c
302e2126
304e20a6
306e2086
1f5c2186
245c005d
345c004e
600c005e
14c36c2c
366441a6
08560496
00000804
f7967016
336460c3
02400f3c
2d72258b
efee103c
080c433c
136414c3
0050313c
313c602e
604e0010
606e6086
3f5c61c6
12c3005d
00c02f3c
343c50c3
61800090
013c00b3
023c013f
23e4016f
780cfb94
06c36c2c
243c15c3
36640090
0e560996
00000804
f8967016
c31750c3
02000f3c
2d72258b
f16e103c
206e2086
1f5c2206
205c0055
305c004e
780c005e
06946047
305c784b
81e6006e
80060173
08946207
6c8c746c
00f00f3c
366416c3
14c383a6
2f3c1364
313c0020
682effc0
ff80313c
740c684e
05c36c2c
24c312c3
08963664
08040e56
fd961016
00c03f3c
4d72458b
fbee233c
4c2e40a6
4c4e4026
4c6e4086
2f5c4266
400c005d
13c3882c
46644126
08560396
00000804
fc961016
326432c3
00076037
60ec2154
04a4335c
1c546007
1a542007
01003f3c
4d72458b
fb6e233c
4c2e40c6
4c4e4046
4c6e4086
2f5c4306
2f5c0075
2f5c0001
400c007d
13c3882c
46644146
001c0073
04960101
08040856
f7961016
0101301c
16540007
02403f3c
4d72458b
efee233c
4c2e40a6
4c4e4026
4c6e4086
2f5c4326
400c005d
13c3882c
46644126
03c330c3
08560996
00000804
f7961016
0101301c
16540007
02403f3c
4d72458b
efee233c
4c2e40a6
4c4e4026
4c6e4086
2f5c43c6
400c005d
13c3882c
46644126
03c330c3
08560996
00000804
fc961016
326432c3
02d26037
001c24f2
03330101
01003f3c
4d72458b
fb6e233c
4c2e40c6
4c4e4046
4c6e40c6
2f5c40a6
2f5c0075
2f5c0001
400c007d
13c3882c
46644146
08560496
00000804
fc961016
326432c3
301c6037
00070101
3f3c1a54
458b0100
233c4d72
40c6fb6e
40464c2e
40c64c4e
41664c6e
00752f5c
00012f5c
007d2f5c
882c400c
414613c3
30c34664
049603c3
08040856
fc963016
201c51c3
00074046
608c1654
121c8c2c
253c00be
3fc30960
20c34664
3f5c0cf2
68120001
00091f5c
155c6c80
31030413
0426355c
049602c3
08040c56
ff963016
4046301c
408c0ed2
0423515c
0ce0313c
880c6037
00ae121c
600625c3
30c34664
019603c3
08040c56
ff963016
4046301c
408c0ed2
0423515c
0ee0313c
880c6037
00ae121c
602625c3
30c34664
019603c3
08040c56
ff961016
4046301c
608c0cd2
0de0213c
8c0c4037
009e121c
60064026
30c34664
019603c3
08040856
ff961016
4046301c
608c0cd2
0be0213c
8c0c4037
009e121c
60064066
30c34664
019603c3
08040856
fe967016
51c340c3
24f202d2
4046001c
604c0a53
121c6c6c
3664009e
4b940007
6c6c704c
153c04c3
36640a60
43940007
6c6c704c
153c04c3
36640ae0
3b940007
6c6c704c
153c04c3
36640b60
33940007
6c6c704c
153c04c3
36640960
2b940007
6fc3704c
04c36c6c
36641fc3
23940007
355c780b
708c0416
04c36c4c
366415c3
19940007
6c6c708c
15c304c3
00073664
708c1294
04c36c8c
366415c3
708c0cf2
04c36cac
366415c3
708c06f2
04c36ccc
366415c3
0e560296
00000804
ff967016
51c360c3
25f202d2
4046201c
0f734037
31c3258b
33647fe5
4d04101c
201c2037
211cfffd
12c30000
6db431e4
604776a9
155c0494
00b30181
21946027
0151155c
341c31c3
60070001
788c1a54
06c36cec
253c15c3
36640ce0
00070037
788c5494
06c38d0c
255c15c3
353c0413
46640960
07f20037
255c4026
00730afd
60376006
604776a9
255c0494
00b30181
21946027
0151255c
341c32c3
60070002
788c1a54
06c36d2c
253c15c3
36640de0
00070037
788c2a94
06c38d4c
3f5c15c3
23c30001
0280363c
00374664
202604f2
0afd155c
604776a9
155c0494
00b30181
13946027
0151155c
341c31c3
6dd20004
6d6c788c
15c306c3
0ee0253c
00373664
402604f2
0afd255c
01960017
08040e56
ff963016
51c340c3
326432c3
001c6037
80070101
345c4454
40062924
0001211c
60073283
70ec1c54
235c4006
70ec0476
235c4006
70ec0447
0484035c
0463135c
08cb9cbc
430670ec
0425235c
50ec702c
023c6c6c
36640440
21940007
15c304c3
00013f5c
78bc23c3
000709bb
345c1894
40062924
0001211c
60073283
702c1054
310c50ec
023c6cac
252c0440
07f23664
235c70ec
43f20473
0444035c
0c560196
00000804
0136f016
50c3fa96
62c381c3
73c36364
305c7364
40062924
0001211c
60073283
60ec1c54
235c4006
60ec0476
235c4006
60ec0447
0484035c
0463135c
08cb9cbc
420674ec
0425235c
54ec742c
023c6c6c
36640440
28940007
00404f3c
231704c3
e6bc4286
803708cb
18c305c3
37c326c3
09bb26bc
18940007
2924355c
211c4006
32830001
10546007
54ec742c
6cac350c
0440023c
3664252c
74ec07f2
0473235c
035c43f2
06960444
0f568076
00000804
40c3f016
52c371c3
636463c3
c4f242d2
0101001c
305c0873
40062924
0001211c
60073283
60ec1c54
235c4006
60ec0476
235c4006
60ec0447
0484035c
0463135c
08cb9cbc
41c670ec
0425235c
50ec702c
023c6c6c
36640440
20940007
17c304c3
36c325c3
09baf4bc
18940007
2924345c
211c4006
32830001
10546007
50ec702c
6cac310c
0440023c
3664252c
70ec07f2
0473235c
035c43f2
0f560444
00000804
40c3f016
62c351c3
73c36364
305c7364
40062924
0001211c
60073283
60ec1c54
235c4006
60ec0476
235c4006
60ec0447
0484035c
0463135c
08cb9cbc
418670ec
0425235c
50ec702c
023c6c6c
36640440
20940007
15c304c3
37c326c3
09bad6bc
18940007
2924345c
211c4006
32830001
10546007
50ec702c
6cac310c
0440023c
3664252c
70ec07f2
0473235c
035c43f2
0f560444
00000804
40c37016
62c351c3
305c6364
40062924
0001211c
60073283
60ec1c54
235c4006
60ec0476
235c4006
60ec0447
0484035c
0463135c
08cb9cbc
414670ec
0425235c
50ec702c
023c6c6c
36640440
1f940007
15c304c3
babc26c3
000709ba
345c1894
40062924
0001211c
60073283
702c1054
310c50ec
023c6cac
252c0440
07f23664
235c70ec
43f20473
0444035c
08040e56
0136f016
50c3fa96
62c381c3
73c36364
305c7364
40062924
0001211c
60073283
60ec1c54
235c4006
60ec0476
235c4006
60ec0447
0484035c
0463135c
08cb9cbc
410674ec
0425235c
54ec742c
023c6c6c
36640440
28940007
00404f3c
231704c3
e6bc4286
803708cb
18c305c3
37c326c3
09ba7abc
18940007
2924355c
211c4006
32830001
10546007
54ec742c
6cac350c
0440023c
3664252c
74ec07f2
0473235c
035c43f2
06960444
0f568076
00000804
40c3f016
62c351c3
73c36364
02d27364
001c24f2
08734046
2924305c
211c4006
32830001
1c546007
400660ec
0476235c
400660ec
0447235c
035c60ec
135c0484
9cbc0463
70ec08cb
235c4086
702c0425
6c6c50ec
0440023c
00073664
04c32094
26c315c3
24bc37c3
000709ba
345c1894
40062924
0001211c
60073283
702c1054
310c50ec
023c6cac
252c0440
07f23664
235c70ec
43f20473
0444035c
08040f56
0336f016
60c3f896
52c371c3
000793c3
20072154
40071f54
60071d54
4f3c1b54
04c30100
9cbc2206
04c308cb
410615c3
08cbb0bc
ac4c784c
17c306c3
3fc324c3
40c35664
09c309f2
42061fc3
08cbb0bc
401c0073
04c34046
c0760896
08040f56
0736f016
60c3f896
af5c81c3
52c30204
93c35364
00079364
20072354
3ac32154
1e546007
20060fc3
bebc4206
4f3c0891
04c30100
9cbc2206
b00e08cb
0016945c
ac4c784c
18c306c3
3fc324c3
40c35664
0ac309f2
42061fc3
08cbb0bc
401c0073
04c34046
e0760896
08040f56
0336f016
50c3f896
72c381c3
9f5c63c3
000701e4
20073254
40073054
60072e54
09c32c54
29540007
01004f3c
220604c3
08cb9cbc
39a26006
602531a1
fc946107
3f3c27c3
023c0180
033c009f
1f3c00df
01c30200
f89430e4
8c4c744c
18c305c3
01002f3c
46643fc3
09f240c3
1fc309c3
b0bc4206
007308cb
4046401c
089604c3
0f56c076
00000804
0336f016
80c3f096
92c361c3
24f202d2
4046401c
0f3c1293
22060300
08cb9cbc
0171065c
141c10c3
20f70001
00612f5c
01852f5c
01c1365c
041c03c3
00b70001
00411f5c
018d1f5c
2f3c56c3
36c30320
03901f3c
0101035c
00df023c
21e46025
4f3cfa94
36c30390
0139135c
00df143c
2f3c6025
02c30400
f79440e4
02000f3c
9cbc2206
165c08cb
1f5c01e1
265c0105
2f5c01e9
365c010d
3f5c01f1
065c0115
0f5c01f9
165c011d
1f5c0201
265c0125
2f5c0209
2f3c012d
36c30260
02c01f3c
0181035c
00df023c
21e46025
3f3cfa94
2c090300
360921c3
40772103
00212f5c
00df233c
34e4a025
18c3f594
7f3c644c
8c4c0100
16c308c3
03002f3c
466437c3
000740c3
50c31c94
02002f3c
03c36aa2
03037ea2
0f5c0037
0aa10001
a207a025
08c3f694
8c4c604c
37c316c3
40c34664
09c306f2
25c317c3
08cbb0bc
109604c3
0f56c076
00000804
0136f016
60c3f796
403771c3
4f3c83c3
04c30140
9cbc2206
04c308cb
40661fc3
08cbb0bc
ac4c784c
17c306c3
3f3c24c3
56640040
2f5c0df2
48120029
00313f5c
69807012
00212f5c
28c36d00
0996680f
0f568076
00000804
f9963016
001c50c3
a0070101
4f3c1c54
658b01c0
343c6d72
62a6f3ee
6226702e
60c6704e
6146706e
005d3f5c
00c00f3c
420612c3
08cbb0bc
6c2c740c
14c305c3
36644326
0c560796
00000804
f996f016
61c350c3
226403c3
a2d24037
001c64f2
05130101
7f3c746c
6ccc0140
366417c3
20940007
01c04f3c
6d72798b
f46e343c
702e6186
704e6106
706e60c6
3f5c6126
3f5c0065
3f5c0001
0f3c006d
17c300e0
b0bc40c6
740c08cb
05c36c2c
420614c3
07963664
08040f56
f9963016
02d250c3
001c44f2
03930101
01c04f3c
6d72658b
f3ee343c
702e62a6
704e6226
706e60c6
3f5c6106
0f3c005d
12c300c0
b0bc4206
740c08cb
05c36c2c
432614c3
07963664
08040c56
fb967016
63c350c3
02d22364
001c64f2
03d30101
01404f3c
6d72658b
f6ee343c
702e61e6
704e6166
706e60c6
3f5c60e6
245c004d
0f3c004e
16c300c0
b0bc4106
740c08cb
05c36c2c
426614c3
05963664
08040e56
f9963016
02d250c3
001c44f2
03730101
01c04f3c
6d72658b
f3ee343c
702e62a6
704e6226
706e60c6
005d3f5c
00c00f3c
420612c3
08cbb0bc
6c2c740c
14c305c3
36644326
0c560796
00000804
f9963016
000750c3
20072154
40071f54
4f3c1d54
658b01c0
343c6d72
62a6f3ee
6226702e
60c6704e
6086706e
005d3f5c
00c00f3c
420612c3
08cbb0bc
6c2c740c
14c305c3
36644326
001c0073
07960101
08040c56
f9963016
000750c3
20072154
40071f54
4f3c1d54
658b01c0
343c6d72
62a6f3ee
6226702e
60c6704e
6066706e
005d3f5c
00c00f3c
420612c3
08cbb0bc
6c2c740c
14c305c3
36644326
001c0073
07960101
08040c56
f9963016
226451c3
326440b7
3f5c6077
60370141
24f202d2
0101401c
2f3c06b3
658b01c0
323c6d72
6166f8ee
60e6682e
60c6684e
6046686e
00ad3f5c
00413f5c
00b53f5c
00213f5c
00bd3f5c
00013f5c
00c53f5c
3f5c6206
315c00cd
3f5c0149
315c00d5
3f5c0151
600c00dd
12c36c2c
366441e6
08f240c3
02b0053c
01501f3c
b0bc40e6
04c308cb
0c560796
00000804
f9963016
226451c3
326440b7
3f5c6077
60370141
24f202d2
0101401c
2f3c0653
658b01c0
323c6d72
6166f8ee
60e6682e
60c6684e
6026686e
00ad3f5c
00413f5c
00b53f5c
00213f5c
00bd3f5c
00013f5c
00c53f5c
3f5c6206
60e600cd
00d53f5c
00dd3f5c
6c2c600c
41e612c3
40c33664
053c08f2
1f3c0240
40e60150
08cbb0bc
079604c3
08040c56
0336f016
71c360c3
92c383c3
4f5c9364
000700e3
00ec4454
04a4305c
3f546007
3d542007
600738c3
80073a54
782c3854
0c856cac
36643fe6
33940007
323c5dab
54c3ffe0
05d434e4
ffd0323c
536453c3
435c78ec
7d8b04a4
700e6d72
0070353c
353c702e
704e0030
706e6086
310d23a6
004e945c
00b0043c
25c318c3
08cbb0bc
6c2c780c
14c306c3
00b0253c
782c3664
6cec58ec
0640023c
00733664
0101001c
0f56c076
00000804
0136f016
40c3ff96
63c381c3
736472c3
00e35f5c
a4f262d2
0101001c
305c08b3
40062924
0001211c
60073283
60ec1c54
235c4006
60ec0476
235c4006
60ec0447
0484035c
0463135c
08cb9cbc
43a670ec
0425235c
50ec702c
023c6c6c
36640440
22940007
00065f5c
18c304c3
36c327c3
09c2ecbc
18940007
2924345c
211c4006
32830001
10546007
50ec702c
6cac310c
0440023c
3664252c
70ec07f2
0473235c
035c43f2
01960444
0f568076
00000804
0336f016
71c360c3
92c383c3
4f5c9364
000700e3
00ec4454
04a4305c
3f546007
3d542007
600738c3
80073a54
782c3854
0c856cac
36643fe6
33940007
323c5dab
54c3ffe0
05d434e4
ffd0323c
536453c3
435c78ec
7d8b04a4
700e6d72
0070353c
353c702e
704e0030
706e6086
310d2366
004e945c
00b0043c
25c318c3
08cbb0bc
6c2c780c
14c306c3
00b0253c
782c3664
6cec58ec
0640023c
00733664
0101001c
0f56c076
00000804
0136f016
81c360c3
000752c3
00ec4954
04a4305c
44546007
42542007
40544007
6cac782c
3fe60c85
00073664
78ec3b94
04a4435c
45ab18c3
323cf44b
37e4ffc0
323c05d4
73c3ffb0
28c37364
6d72698b
344b700e
612531c3
544b702e
60a532c3
6086704e
22e6706e
540b310d
004e245c
345c742b
043c005e
344c00d0
b0bc27c3
780c08cb
06c36c2c
273c14c3
366400d0
58ec782c
023c6cec
36640640
001c0073
80760101
08040f56
0136f016
81c350c3
000772c3
00ec4754
04a4305c
42546007
40542007
3e544007
6cac742c
3fe60c85
00073664
18c33994
dc4b45ab
ffc0323c
05d436e4
ffb0323c
636463c3
435c74ec
28c304a4
6d72698b
363c700e
702e0090
0050363c
6086704e
22c6706e
5c0b310d
004e245c
345c7c2b
043c005e
3c4c00d0
b0bc26c3
740c08cb
05c36c2c
263c14c3
366400d0
54ec742c
023c6cec
36640640
001c0073
80760101
08040f56
40c37016
62c351c3
44f222d2
0101001c
305c0853
40062924
0001211c
60073283
60ec1c54
235c4006
60ec0476
235c4006
60ec0447
0484035c
0463135c
08cb9cbc
42c670ec
0425235c
50ec702c
023c6c6c
36640440
1f940007
15c304c3
40bc26c3
000709c4
345c1894
40062924
0001211c
60073283
702c1054
310c50ec
023c6cac
252c0440
07f23664
235c70ec
43f20473
0444035c
08040e56
0336f016
71c360c3
92c383c3
4f5c9364
000700e3
00ec4254
04a4305c
3d546007
3b542007
600738c3
782c3854
0c856cac
36643fe6
33940007
323c5dab
54c3ffe0
05d434e4
ffd0323c
536453c3
435c78ec
7d8b04a4
700e6d72
0070353c
353c702e
704e0030
706e6086
310d2a46
004e945c
00b0043c
25c318c3
08cbb0bc
6c2c780c
14c306c3
00b0253c
782c3664
6cec58ec
0640023c
00733664
0101001c
0f56c076
00000804
0336f016
71c360c3
92c383c3
5f5c9364
000700e3
00ec4254
04a4305c
3d546007
3b542007
600738c3
782c3854
0c856cac
36643fe6
33940007
435c78ec
5dab04a4
ffe0323c
05d435e4
ffd0323c
536453c3
6d727d8b
353c700e
702e0070
0030353c
6086704e
2246706e
945c310d
043c004e
18c300b0
b0bc25c3
780c08cb
00b0253c
06c36c2c
236414c3
782c3664
6cec58ec
0640023c
00733664
0101001c
0f56c076
00000804
0136f016
40c3ff96
63c381c3
736472c3
00e35f5c
a4f262d2
0101001c
305c08b3
40062924
0001211c
60073283
60ec1c54
235c4006
60ec0476
235c4006
60ec0447
0484035c
0463135c
08cb9cbc
424670ec
0425235c
50ec702c
023c6c6c
36640440
22940007
00065f5c
18c304c3
36c327c3
09c530bc
18940007
2924345c
211c4006
32830001
10546007
50ec702c
6cac310c
0440023c
3664252c
70ec07f2
0473235c
035c43f2
01960444
0f568076
00000804
0136f016
60c3ff96
83c371c3
40372264
00e14f5c
45540007
305c00ec
600704a4
20074054
18c33e54
3b542007
39548007
6cac782c
3fe60c85
00073664
5dab3494
fff0323c
34e454c3
323c05d4
53c3ffe0
78ec5364
04a4435c
6d727d8b
353c700e
702e0060
0020353c
6086704e
2226706e
3f5c310d
712d0001
00a0043c
25c318c3
08cbb0bc
6c2c780c
14c306c3
00a0253c
782c3664
6cec58ec
0640023c
00733664
0101001c
80760196
08040f56
0136f016
50c3ff96
82c371c3
236423c3
40540007
305c00ec
600704a4
20073b54
18c33954
36542007
34544007
6cac742c
3fe60c85
36644037
00074017
7dab2d94
32e462c3
7fe504d4
636463c3
435c74ec
7d8b04a4
700e6d72
0050363c
363c702e
704e0010
706e6086
310d21e6
0090043c
b0bc18c3
740c08cb
05c36c2c
263c14c3
36640090
54ec742c
023c6cec
36640640
001c0073
01960101
0f568076
00000804
0136f016
50c3fe96
82c371c3
60773364
44540007
305c00ec
600704a4
20073f54
40073d54
20573b54
38542007
6cac742c
3fe60c85
00073664
7dab3394
00216f5c
12c34057
06d431e4
fff0133c
6f5c2037
74ec0001
04a4435c
6d727d8b
363c700e
702e0050
0010363c
4086704e
61a6506e
043c710d
18c30090
b0bc26c3
740c08cb
05c36c2c
263c14c3
36640090
54ec742c
023c6cec
36640640
001c0073
02960101
0f568076
00000804
0136f016
71c360c3
53c382c3
00075364
00ec3d54
04a4305c
38546007
36542007
34544007
3254a007
6cac782c
3fe60c85
00073664
78ec2d94
04a4435c
35e47dab
7fe504d4
536453c3
6d727d8b
353c700e
702e0050
0010353c
6086704e
4166706e
043c510d
18c30090
b0bc25c3
780c08cb
06c36c2c
253c14c3
36640090
58ec782c
023c6cec
36640640
001c0073
80760101
08040f56
0136f016
60c3ff96
83c371c3
226481d7
00074037
00ec4254
04a4305c
3d546007
3b542007
400728c3
80073854
782c3654
0c856cac
36643fe6
31940007
535c78ec
5dab04a4
7fc532c3
023543e4
436443c3
6d727d8b
343c740e
742e0060
0020343c
6086744e
4126746e
3f5c550d
752d0001
00a0053c
24c318c3
08cbb0bc
6c2c780c
15c306c3
00a0243c
782c3664
6cec58ec
0640023c
00733664
0101001c
80760196
08040f56
f8967016
01c360c3
c00712c3
00073754
40073554
41ab3354
323ca46b
35e4ffa0
323c05d4
53c3ff90
4f3c5364
618b0200
343c6d72
646bf0ee
00b0233c
60e5502e
6086704e
60c6706e
004d3f5c
345c640b
642b004e
005e345c
345c644b
0f3c006e
244c0100
b0bc25c3
780c08cb
06c36c2c
253c14c3
366400f0
001c0073
08960101
08040e56
40c37016
62c351c3
45540007
43542007
41544007
2924305c
211c4006
32830001
1c546007
400660ec
0476235c
400660ec
0447235c
035c60ec
135c0484
9cbc0463
70ec08cb
235c40c6
702c0425
6c6c50ec
0440023c
00073664
04c32094
26c315c3
09c770bc
2924345c
211c4006
32830001
13546007
50ec702c
6cac310c
0440023c
3664252c
70ec0af2
0473235c
035c46f2
00730444
0101001c
08040e56
0136f016
60c3ff96
83c371c3
40372264
00e35f5c
44540007
305c00ec
600704a4
20073f54
18c33d54
3a542007
3854a007
6cac782c
3fe60c85
00073664
78ec3394
04a4435c
323c5dab
35e4fff0
323c05d4
53c3ffe0
7d8b5364
700e6d72
0060353c
353c702e
704e0020
706e6086
310d20a6
00013f5c
043c712d
18c300a0
b0bc25c3
780c08cb
06c36c2c
253c14c3
366400a0
58ec782c
023c6cec
36640640
001c0073
01960101
0f568076
00000804
50c33016
013c41c3
15c30100
b0bc4086
043c08cb
153c00e0
40460040
08cbb0bc
00c0043c
0060153c
b0bc4046
043c08cb
153c00a0
40460080
08cbb0bc
0080043c
00a0153c
b0bc4046
043c08cb
153c0040
408600c0
08cbb0bc
0c560006
00000804
50c33016
220541c3
b0bc4086
053c08cb
143c0040
404600e0
08cbb0bc
0060053c
00c0143c
b0bc4046
053c08cb
143c0080
404600a0
08cbb0bc
00a0053c
0080143c
b0bc4046
053c08cb
143c00c0
40860040
08cbb0bc
0c560006
00000804
1f36f016
90c3f496
00ec71c3
501c80b0
20074046
606c4754
21456c4c
60c33664
4d05501c
3e540007
4d04501c
2007218b
2cc33954
39c30870
b75cacec
a75c0033
20460043
201c21f7
2f5c2800
4f3c0106
04c30080
01c01f3c
e6bc4286
803708cb
16c305c3
3ac32bc3
50c38664
0cec39c3
2924305c
111c2006
31830001
12546007
1094a007
7c8940ec
85cc1cc3
0484025c
0473125c
46645c0c
00770364
00212f5c
05c35cad
f8760c96
08040f56
f5967016
41c360c3
24f202d2
4046001c
60ec09b3
484c4c6c
210503c3
50c32664
4d05001c
4254a007
4d04001c
2007358b
500b3d54
01062f5c
3f5c702b
101c0116
1f5c2800
302c0126
2f5c444b
0f3c0136
02b70020
6047642c
648b0494
0113600e
06946207
6c6c78ec
20856c8c
58ec3664
6c2c68ac
15c302c3
02002f3c
38ec3664
2924315c
211c4006
32830001
0ef26fd2
64ec502c
0484335c
280e2c0b
78ec502c
335c6cec
2c2b0484
0b96282e
08040e56
1f36f016
90c3f596
00ec71c3
501c80b0
20074046
606c4154
21856c4c
60c33664
4d05501c
38540007
4d04501c
4007418b
3cc33354
29c30c50
b75ca8ec
a75c0003
60460013
201c61b7
2f5c2802
4f3c00e6
04c30040
01801f3c
e6bc4286
803708cb
16c305c3
3ac32bc3
50c38664
0cec39c3
2924305c
211c4006
32830001
acf26dd2
2cc360ec
035c89ec
135c0484
5c2c0473
46647c8b
05c31cae
f8760b96
08040f56
1f36f016
90c3f596
00ec71c3
501c80b0
20074046
606c4154
21856c4c
60c33664
4d05501c
38540007
4d04501c
4007418b
3cc33354
29c30c50
b75ca8ec
a75c0003
60460013
201c61b7
2f5c2803
4f3c00e6
04c30040
01801f3c
e6bc4286
803708cb
16c305c3
3ac32bc3
50c38664
0cec39c3
2924305c
211c4006
32830001
acf26dd2
2cc360ec
035c8a0c
135c0484
5c2c0473
46647c8b
05c31cae
f8760b96
08040f56
0136f016
51c370c3
00b000ec
4046601c
2a542007
6c4c606c
36642185
601c10c3
00074d05
601c2154
418b4d04
1c544007
8c0c38c3
540b1cec
4664742b
1cec60c3
2924305c
211c4006
32830001
ccf26dd2
28c360ec
035c8a2c
135c0484
542c0473
4664748b
06c314ae
0f568076
00000804
ff967016
41c350c3
24f202d2
4046001c
60ec0393
484c4c6c
214503c3
10c32664
4d05001c
11542007
4d04001c
6dd2658b
4cac74ec
d02cb00b
0f5c108b
890c0006
25c303c3
466436c3
0e560196
00000804
ff967016
41c350c3
24f202d2
4046001c
60ec0393
484c4c6c
214503c3
10c32664
4d05001c
11542007
4d04001c
6dd2658b
4cac74ec
d02cb00b
0f5c108b
892c0006
25c303c3
466436c3
0e560196
00000804
0336f016
70c3fd96
02d241c3
001c24f2
08534046
4c6c60ec
03c3484c
26642145
600650c3
4d05001c
2794a007
49a006b3
21e42246
12c303d4
558b1164
2a544007
0f5c100b
83c30006
08c38364
6100502b
00163f5c
636461c3
00266f5c
60b7702c
68ac5cec
02c36d4c
2fc315c3
00073664
08c31394
31647800
32e4508b
558bd974
7cec49d2
896c4cac
15c303c3
46644026
001c0073
03964d04
0f56c076
00000804
ff967016
41c350c3
24f202d2
4046001c
60ec0393
484c4c6c
214503c3
10c32664
4d05001c
11542007
4d04001c
6dd2658b
4cac74ec
d02cb00b
0f5c108b
898c0006
25c303c3
466436c3
0e560196
00000804
ff967016
41c350c3
24f202d2
4046001c
60ec0393
484c4c6c
214503c3
10c32664
4d05001c
11542007
4d04001c
6dd2658b
4cac74ec
d02cb00b
0f5c108b
89ac0006
25c303c3
466436c3
0e560196
00000804
60c3f016
02d251c3
401c24f2
07934046
4c6c60ec
03c3484c
26642285
401c10c3
00074d05
401c3154
618b4d04
2c546007
f52ee006
68ac58ec
02c38cec
74ab25c3
40c34664
325c58ec
20062924
0001111c
60073183
00071954
68ec1794
0473035c
21c3350b
30c32364
23e43364
10c30235
236421c3
48d2552e
6cec78ec
135c146c
b0bc0484
04c308cb
08040f56
60c3f016
02d251c3
401c24f2
07534046
4c6c60ec
03c3484c
26642185
401c10c3
00074d05
401c2f54
618b4d04
2a546007
68ac58ec
02c38ccc
74ab540b
40c34664
325c58ec
e0062924
0001711c
60073783
00071954
68ec1794
0473035c
21c3348b
30c32364
23e43364
10c30235
336431c3
58ec74ae
142c48ec
0484125c
b0bc23c3
04c308cb
08040f56
60c3f016
02d251c3
401c24f2
07334046
4c6c60ec
03c3484c
26642185
401c10c3
00074d05
401c2e54
618b4d04
29546007
68ac58ec
02c36c8c
3664540b
58ec40c3
2924325c
711ce006
37830001
19546007
17940007
035c68ec
348b0473
236421c3
336430c3
023523e4
31c310c3
74ae3364
48ec58ec
125c142c
23c30484
08cbb0bc
0f5604c3
00000804
0336f016
50c3fa96
02d271c3
401c24f2
09534046
4c6c60ec
03c3484c
26642405
401c60c3
00074d05
401c3f54
218b4d04
3a542007
4f3c14f0
04c30040
0040173c
e6bc4286
28c308cb
5c0b68ac
0013975c
8c4c8037
16c308c3
466439c3
54ec40c3
2924325c
611cc006
36830001
1c546007
1a940007
335c68ec
6c090484
1dcb13c3
236423c3
336430c3
023523e4
21c310c3
5dee2364
6cec74ec
0484335c
133c1ccc
b0bc0010
04c308cb
c0760696
08040f56
0736f016
70c3fd96
a364a1c3
936493c3
0001805c
c00652c3
05738026
540e5e62
0020043c
4f5c00b7
831c0041
0a940001
542f4046
748e7e62
20773100
00214f5c
831c0233
0e940002
020635c3
027e033c
13c31e00
09c856bc
0100243c
4f5c4037
363c0001
63c30010
a3056364
053469e4
336434c3
d3143ae4
039606c3
0f56e076
00000804
0736f016
60c3fb96
a364a1c3
936493c3
0001805c
802652c3
0733e006
540e5a62
0020043c
3f5c0137
39a20081
033c348d
00f70010
00613f5c
346e39e2
0020033c
4f5c00b7
831c0041
0a940007
544f4046
74ce7a62
20773100
00214f5c
831c0233
0e940015
020635c3
047e033c
13c31a00
09c856bc
0100243c
4f5c4037
373c0001
73c30010
a3857364
053479e4
336434c3
c5143ae4
059607c3
0f56e076
00000804
0736f016
a1c360c3
93c3a364
805c9364
52c30001
8026e006
5a620553
343c540e
33640020
142e19e2
43c36045
831c4364
07940006
542f4046
748e7a62
01d37100
0014831c
35c30d94
133c2206
1a00027e
56bc13c3
343c09c8
43c30100
373c4364
73c30010
a3057364
033479e4
d6144ae4
e07607c3
08040f56
0736f016
60c3fb96
a364a1c3
936493c3
0001805c
802652c3
0893e006
540e5a62
0020043c
3f5c0137
39e20081
033c344e
00f70020
00613f5c
346e39e2
0020033c
4f5c00b7
831c0041
09940006
544f4006
00c0053c
9cbc2206
03b308cb
0008831c
00460a94
3a62144f
700034ce
4f5c6077
02330021
0016831c
35c30e94
133c2206
1a00047e
56bc13c3
343c09c8
60370100
00014f5c
0010373c
736473c3
79e4a385
34c30534
3ae43364
07c3ba14
e0760596
08040f56
24f202d2
4046001c
60cc0233
20cf69f2
458b20ef
458b420e
03c3422e
60ec00f3
20ef2d8f
622e658b
08040006
0136f016
60c3ff96
53c381c3
736472c3
34542007
32540007
30546007
6ccc60cc
36641fc3
03f240c3
05530017
602d6046
6046e18e
301c60ef
620e2802
740b20c3
016e323c
682e742b
6086342c
20472ed2
748b0594
60c6684e
786c0113
00c56c8c
0040153c
62863664
6006716e
78cc718f
08c36c2c
366414c3
001c0073
01964046
0f568076
00000804
0136f016
60c3ff96
53c381c3
736472c3
37542007
35540007
33546007
6ccc60cc
36641fc3
03f240c3
05b30017
202d2046
4046e18e
301c40ef
620e2803
340930c3
015e133c
235c542b
542c000e
06944047
235c548b
60a6001e
60660173
08944207
6c8c786c
153c00a5
36640040
716e6266
518f4006
6c2c78cc
14c308c3
00733664
4046001c
80760196
08040f56
0136f016
70c3f996
83c342c3
536451c3
680c03d2
201c66f2
18c34046
0873440f
6c8c60cc
366418c3
000760c3
531c3d54
1c942800
00805f3c
14c305c3
e6bc4286
7ccc08cb
07c38c4c
5a2b16c3
466435c3
040f18c3
27940007
4c097d0c
202512c3
2f5c2077
4c0d0021
531c03f3
1c942801
00805f3c
14c305c3
e6bc4286
7ccc08cb
07c38c6c
5a2b16c3
466435c3
040f18c3
7d0c0af2
12c34c29
20372025
00012f5c
00534c2d
06c3c006
80760796
08040f56
41c31016
60cc4364
14c36c0c
20c33664
40cc07d2
34e4698b
498c0354
02c35cf2
08040856
60ccff96
36646cac
13540007
32c34029
0010341c
018c6ed2
620b0cd2
2902331c
60060894
002b6037
05940027
00730037
60376006
00012f5c
019602c3
00000804
60ccff96
36646cac
12540007
31c32029
0020341c
018c6dd2
620b0bd2
2902331c
602b0794
233c6132
40370014
60060073
1f5c6037
01c30001
08040196
842b7016
c42ca48b
48ac40cc
2664240b
001c30c3
60074d06
4d6b1354
42e44fd2
4a200db4
0ad425e4
033c6e00
16c30020
b0bc2364
000608cb
001c0073
0e564046
00000804
41c33016
6cac60cc
3664240b
001c50c3
a0074d06
556b1754
12544007
12e4302b
48a00fb4
23e4708b
23640bd4
748050ae
133c102c
b0bc0020
000608cb
001c0073
0c564046
00000804
0736f016
60c3fe96
32c3a1c3
40374909
0003835c
ac6cec2c
0083935c
04f222d2
4046001c
60cc0553
1f3c6ccc
36640040
03f240c3
04330057
00013f5c
805c602d
37c300c6
024f233c
040540ef
420613c3
08cbb0bc
043caad2
15c30020
b0bc29c3
945c08cb
005300b6
6006b16e
78cc718f
0ac36c2c
366414c3
e0760296
08040f56
0136f016
70c3ff96
63c381c3
536452c3
38540007
36542007
60076c0c
60cc3354
1fc36ccc
40c33664
001703f2
404605b3
a18e402d
60ef6046
2801201c
083c420e
16c30040
b0bc4286
404608cb
4c2d38c3
a047b80c
584b0494
0153502e
a2076006
7c6c0894
043c6c8c
16c30020
35c33664
6006716e
7ccc718f
08c36c2c
366414c3
001c0073
01964046
0f568076
00000804
0136f016
70c3ff96
63c381c3
536452c3
38542007
36540007
60076c0c
60cc3354
1fc36ccc
40c33664
001703f2
404605b3
a18e402d
60ef6046
2800201c
083c420e
16c30040
b0bc4286
402608cb
4c2d38c3
a047b80c
584b0494
0153502e
a2076006
7c6c0894
043c6c8c
16c30020
35c33664
6006716e
7ccc718f
08c36c2c
366414c3
001c0073
01964046
0f568076
00000804
fa96f016
71c360c3
24f202d2
4046001c
406c0c33
bc0b2449
01403f3c
880c6037
0030273c
466435c3
000750c3
784c1394
06c36c2c
42663c0b
18ec3664
323c4289
66d20044
41374292
00811f5c
0157228d
403c0833
04c30420
9cbc2206
784c08cb
06c36c6c
366414c3
34940007
784c0177
06c36c6c
04a0153c
00073664
01772b94
4e8978ec
341c32c3
6cd20004
76ad6046
2e8978ec
241c21c3
40f700fb
00611f5c
78ec2e8d
32c34e89
0001341c
60266cd2
78ec76ad
21c32e89
00fe241c
1f5c40b7
2e8d0041
4e8978ec
40774372
00211f5c
06962e8d
08040f56
17df83ff
d14e0932
918acde7
c4c4d5c6
4e182140
dcf48655
eca7158a
5393df92
34ca1830
59c7a2bf
0dba8f67
7d2dd86d
97570a54
7ad23970
853324ea
e11d9aed
2ebe07ff
a39d1264
23159bcf
8889ab8d
9c304280
b9e90dab
d94f2b14
a626bf25
69943160
b28e457f
1a741fcf
fa5ab0db
2eaf14a8
f5a473e0
0b6748d4
c33b34db
5c7c0ffe
473b25c8
472a369f
1113571b
39618400
72d31b56
b29f5628
4c4d7e4b
d22863c0
651d8bfe
35e83e9e
f5b560b7
5d5e2950
eb49e7c0
17ce90a8
877768b6
b9f81efc
8f764a90
8e546c3e
2226ae36
72c20801
e4a637ac
643fad50
999afc96
a551c680
cb3a16fd
6bd07d3c
ea6bc16e
bbbc52a0
d793ce81
2f9c2151
00efd06c
0400feff
50001800
4004e001
01558019
180404fe
e1515018
995944e4
faff54d5
48001c00
a005b001
814cc01d
1cfa05ab
b149481c
ddbda5b5
ae2acd8c
5400e6ff
1004f801
41516018
195184e7
f95554e6
780814fc
63a61031
b2ff48d5
e805ac01
2149701c
9db6c5b6
adb34db7
6cf4eda9
73976839
fa2a2b73
44041efe
51559819
5800e4ff
e004d001
815d401a
1bae04cd
d15958e4
5afae4d4
c94cdc1d
bcffb5aa
30058801
c147a01e
1f638590
89bd434a
be2e358d
155186e7
09557ce6
b80434fe
6159901b
9af344d7
caf75c29
8ba3bc30
93b638c9
75b369b7
8cfa3dab
f142281f
de24258e
96dec6da
379376c7
ab7fb36a
1c04fa01
b1514818
d95da4e5
00aad4cc
e8fbc1ff
8b72904c
8951b3e7
2323ab63
72188402
3b2f61aa
37e5a851
cac9fb49
2c53180c
9ae345fd
b05df1e6
beb41bb6
e9ea502a
5e4b9c0e
a1cc2457
87b859b7
747de0ff
c5b94826
c4a8d9f3
1191d5b1
390c4201
9d97b0d5
9bf2d428
6564fda4
96298c06
4d71a2fe
582ef8f3
5f5a0ddb
74f52815
af25ce07
d0e6122b
c3dc2cdb
3a3ef07f
e2dca413
e2546cf9
88c8ead8
9c862100
4ecbd86a
4df96a14
32b27ed2
4b14c603
a6b8d17f
ac177c79
afad06ed
ba7a940a
d792e703
e8730915
e1ee166d
9d1f783f
f16e5209
712a367c
4464756c
4e431080
2765ec35
26fcb50a
99593f69
a58a6301
d35c68bf
d60bbe3c
57d68376
dd3d4a05
ebc97381
f439848a
f0f70b36
ce8fbc1f
78b72904
38951b3e
22323ab6
a7218840
13b2f61a
937e5a85
ccac9fb4
d2c53180
69ae345f
6b05df1e
abeb41bb
ee9ea502
75e4b9c0
7a1cc245
f87b859b
6747de0f
3c5b9482
1c4a8d9f
11191d5b
5390c420
89d97b0d
49bf2d42
66564fda
e96298c0
34d71a2f
b582ef8f
55f5a0dd
774f5281
baf25ce0
bd0e6122
fc3dc2cd
33a3ef07
9e2dca41
8e2546cf
088c8ead
a9c86210
44ecbd86
24df96a1
332b27ed
f4b14c60
9a6b8d17
dac177c7
aafad06e
3ba7a940
5d792e70
de873091
fe1ee166
99d1f783
cf16e520
c712a367
04464756
54e43108
a2765ec3
926fcb50
199593f6
fa58a630
cd35c68b
6d60bbe3
557d6837
1dd3d4a0
aebc9738
6f439848
ff0f70b3
4ce8fbc1
e78b7290
638951b3
022323ab
aa721884
513b2f61
4937e5a8
0ccac9fb
fd2c5318
e69ae345
b6b05df1
2abeb41b
0ee9ea50
575e4b9c
b7a1cc24
ff87b859
26747de0
f3c5b948
b1c4a8d9
011191d5
d5390c42
289d97b0
a49bf2d4
066564fd
fe96298c
f34d71a2
db582ef8
155f5a0d
0774f528
2baf25ce
dbd0e612
7fc3dc2c
133a3ef0
f9e2dca4
d8e2546c
0088c8ea
6a9c8621
144ecbd8
d24df96a
0332b27e
7f4b14c6
79a6b8d1
edac177c
0aafad06
03ba7a94
15d792e7
6de87309
3fe1ee16
099d1f78
7cf16e52
6c712a36
80446475
354e4310
0a2765ec
6926fcb5
0199593f
bfa58a63
3cd35c68
76d60bbe
0557d683
81dd3d4a
8aebc973
36f43984
1ff0f70b
04ce8fbc
3e78b729
b638951b
4022323a
1aa72188
8513b2f6
b4937e5a
80ccac9f
5fd2c531
1e69ae34
bb6b05df
02abeb41
c0ee9ea5
4575e4b9
9b7a1cc2
0ff87b85
826747de
9f3c5b94
5b1c4a8d
2011191d
0d5390c4
4289d97b
da49bf2d
c066564f
2fe96298
8f34d71a
ddb582ef
8155f5a0
e0774f52
22baf25c
cdbd0e61
07fc3dc2
4133a3ef
cf9e2dca
ad8e2546
10088c8e
86a9c862
a144ecbd
ed24df96
60332b27
17f4b14c
c79a6b8d
6edac177
40aafad0
703ba7a9
915d792e
66de8730
83fe1ee1
2099d1f7
67cf16e5
56c712a3
08044647
c354e431
50a2765e
f6926fcb
30199593
8bfa58a6
e3cd35c6
376d60bb
a0557d68
381dd3d4
48aebc97
b36f4398
00000070
0013a978
93e22d01
ae1545be
a4870378
3fcf38b8
94096708
6ba826eb
1b3418bd
f772bfbb
9c483540
553b2f51
d89fc0e3
b18df3d3
dc3ea7ff
a6d77786
baf4fb11
83649192
daef33f1
2bb2b52c
cb99d188
141d848c
ca719781
578ba35f
52c4823c
a0e81c5c
4a85b404
b65413f6
8e1a0cdf
fc39e0de
4e249b20
ab9e98a9
6cd060f2
d9c7faea
6e1fd400
53ecbc43
5d7afe89
c232c949
6df89af9
9659db16
e6cde944
0a8f4246
65b9ccc1
acc6d2b0
2962411e
50740e2e
25c35a02
5b2a8a7b
470d06f0
7e9d706f
2712ce10
d64f4cd5
36683079
ede47d75
37906a80
aa765ea2
af3d7fc5
6119e5a5
b77c4dfd
4badee0b
73e7f522
05c82123
b3dd66e1
56636958
9531a10f
283a0717
09b00080
fdb9ef60
e49f1210
f8adba69
65c238c0
fc94064f
1b6ade19
82a84e5d
ece8ed70
c315b372
47b6abff
25ac0144
418efac9
d3cb211a
26fe6e0d
0f32da58
849da920
bb9c0598
e7638c22
c673e1c5
875b24af
57f72766
b7b196f4
54d58b5c
f6aadf79
11f1a33e
17d1f5ca
bc83937b
eb1e52bd
35d6ccae
b48ac808
d9bfcde2
3f5950d0
0a34624d
56b58848
9e6b2e4c
033c3dd2
5197fb13
71914a75
2a76be23
55d4f95f
3137dc0b
77d77416
db07e6a7
f3462fa4
e3674561
1c3ba20c
1d041885
b28fa029
7ea6d85a
4b538dee
0ec19aa1
2ca5497a
36c7c481
95437f2b
686cf233
2802f06d
ea9bddce
147c995e
42e5cf86
2d7840b8
1f64e93a
397d9092
3089e06f
bab19746
0a10b7a3
c9b337c5
64ac285a
c6aaabec
0d589567
6ef69af8
3d05dc66
89d8c38a
4936e96a
d4ebbf43
a0689b96
1f92575d
bb5c71d5
7bbec122
946399bc
34b8612a
fbfd1932
51e64017
8f44411d
de8004dd
7fd631e7
39f7a201
ca236fda
d11cd03a
a1123e30
a8e00fcd
2c5982af
efb2ad7d
75ce87c2
90021306
33722e4f
a9cf8dc0
27c4e281
9f7a6c2f
3815e152
c74220fc
5509e408
76148c5e
d7dfff60
00210bfa
b9a6f91a
4c629ee8
d25091d9
8407b418
c8a45bea
6948cb0e
359c4e4b
e5544d45
4a0c3c25
a7cc3f8b
f4ae6bdb
6d7cf32d
7426b59d
b05393f2
83ed11f0
731603b6
708e1e3b
471b86bd
f156247e
b1974688
10b7a3ba
b337c50a
ac285ac9
6a09e667
bb67ae85
3c6ef372
a54ff53a
510e527f
9b05688c
1f83d9ab
5be0cd19
428a2f98
71374491
b5c0fbcf
e9b5dba5
3956c25b
59f111f1
923f82a4
ab1c5ed5
d807aa98
12835b01
243185be
550c7dc3
72be5d74
80deb1fe
9bdc06a7
c19bf174
e49b69c1
efbe4786
0fc19dc6
240ca1cc
2de92c6f
4a7484aa
5cb0a9dc
76f988da
983e5152
a831c66d
b00327c8
bf597fc7
c6e00bf3
d5a79147
06ca6351
14292967
27b70a85
2e1b2138
4d2c6dfc
53380d13
650a7354
766a0abb
81c2c92e
92722c85
a2bfe8a1
a81a664b
c24b8b70
c76c51a3
d192e819
d6990624
f40e3585
106aa070
19a4c116
1e376c08
2748774c
34b0bcb5
391c0cb3
4ed8aa4a
5b9cca4f
682e6ff3
748f82ee
78a5636f
84c87814
8cc70208
90befffa
a4506ceb
bef9a3f7
c67178f2
52c37016
f524ce24
6cd2604c
604f7fe5
233c608c
440f0040
408f4c0c
40060c0f
420606b3
3254a007
11b4301c
0000311c
301c8c0c
311cab40
734f0013
33ef136f
323c412c
612f0010
810f45f2
93af938f
610c00f3
4fac738f
8b8f53af
41068faf
6026518f
b26f71cf
1250201c
0000211c
6025680c
363c680f
62d24004
04c3f324
09f1a4bc
0424245c
363c00b3
62d24004
02c3f324
08040e56
436c3016
36544007
f5248e24
6007634c
680c2d54
4f43101c
424c111c
35e451c3
20062594
692c234f
692f7fe5
690f63f2
238c0133
67af63ac
690c2f8f
029430e4
618c290f
12946107
205c4206
201c0427
211c1250
680c0000
680f6025
4004343c
f32462d2
09f102bc
343c00b3
62d24004
0c56f324
00000804
0136f016
51c360c3
73c342c3
46062006
0891b0bc
5f868065
61974283
b82f3283
78cff8af
043c98ef
141d0040
5c005300
200637c3
202500b3
32c34c0f
15e44800
6e20fb14
235c4006
b84fffe7
00a6b86f
2654a007
0e24f88f
301cf524
311c4f43
780f424c
11a4301c
0000311c
213c2c0c
4c0f0010
11a0301c
0000311c
cc0f25f2
d96fd94f
6c0c00f3
cd6f4d6c
596fc94f
303c794f
03c34004
f32463d2
80760006
08040f56
ae24f016
6006f524
201c600f
211c11a4
680c0000
680f7fe5
11a0101c
0000111c
640f63f2
414c0133
696f616c
640c4d4f
029430e4
201c440f
211c1250
680c0000
680f6025
6006410c
812c610f
353c612f
60074004
f3241554
f5240273
6b4f6006
325c6026
ab8c0427
60257c0c
c2d27c0f
02c3f324
09f102bc
25c39fe5
701c0113
711c1250
6e240000
4004633c
1250101c
0000111c
e2948007
f5244e24
7fe5640c
323c640f
62d24004
e4bcf324
000609f0
08040f56
0136f016
c1d7a197
8e24e217
f52484c3
802c23d2
43d2840f
280f204c
406c63d2
a3d24c0f
740f610c
812cc3d2
e3d2980f
3c0f214c
4004383c
f32462d2
80760006
08040f56
00000804
0736f016
ce2450c3
e12cf524
07b4e027
4004363c
53546007
0a33f324
e047550c
2b8c0e94
896c656c
39e494c3
350f0234
4004363c
43546007
0833f324
0b8c42c3
1250301c
0000311c
40254c0c
550c4c0f
86c314c3
656c4170
a9e493c3
10c30234
4004363c
f32462d2
f52468c3
079442e4
94c3952c
039479e4
0093038c
0b8cf52c
02e412c3
42c30354
301cfcd3
311c1250
4c0c0000
4c0f5fe5
0b5410e4
47ac678c
6b8f4faf
078f63ac
2f8f67af
350f23af
4004383c
f32462d2
09f0e4bc
e0760006
08040f56
10c31016
f5248e24
233c30c3
090cfe4e
21540007
7fe5692c
63f2692f
00d3690f
690f638c
4faf43ac
60066b8f
63ec634f
20062c0f
0427105c
1250201c
0000211c
6025680c
343c680f
62d24004
02bcf324
017309f1
2c0f288c
684c688f
684f6025
4004343c
f32462d2
08560006
00000804
40c33016
25540007
001c600c
011c4f43
50c3424c
1d9435e4
20070066
40071d54
301c1454
311c139c
6c0c0000
13946007
11b4301c
0000311c
001c6c0c
011c12c0
50c30000
075435e4
54bc04c3
009309d5
00530046
0c560086
00000804
0336f016
50c3ff96
62c381c3
9f5c73c3
00070104
62576554
62946607
f5242e24
1250201c
0000211c
6025680c
313c680f
62d24004
301cf324
311c11a0
8c0c0000
11a4301c
0000311c
40066c0c
54e400b3
914c0554
23e44025
2e24fb14
201cf524
211c1250
680c0000
680f7fe5
4004313c
f32462d2
09f0e4bc
325454e4
e0070066
36c33254
31833f86
0040233c
3f8639c3
00a63183
27b423e4
11b4301c
0000311c
201c6c0c
211c12c0
12c30000
1a5431e4
139c201c
0000211c
69d2680c
201c680c
211cf0ef
12c3f0f0
0c3531e4
00079f5c
18c305c3
37c326c3
09d5dcbc
00460093
02660053
c0760196
08040f56
1f540007
101c600c
111c4f43
21c3424c
179432e4
139c301c
0000311c
60076c0c
301c1294
311c11b4
6c0c0000
12c0101c
0000111c
32e421c3
2ebc0654
009309d6
00530046
08040266
fd967016
12540007
501c800c
511c4f43
65c3424c
0a9446e4
803781d7
a077a217
c0b7c257
09d688bc
00460053
0e560396
00000804
600c0cd2
4f43101c
424c111c
32e421c3
acbc0494
005309d6
08040046
305c0fd2
6cd2ffe4
101c6c0c
111c4f43
21c3424c
049432e4
09d70ebc
00660053
00000804
50c37016
000761c3
45075254
2e245094
201cf524
211c1250
680c0000
680f6025
4004313c
f32462d2
1190301c
0000311c
301c8c0c
311c1194
6c0c0000
00b34006
055454e4
402590cc
fb1423e4
f5242e24
1250201c
0000211c
7fe5680c
313c680f
62d24004
e4bcf324
54e409f0
301c2054
311c11b4
6c0c0000
12c0101c
0000111c
32e421c3
201c1654
211c139c
680c0000
680c69d2
f0ef101c
f0f0111c
32e421c3
05c30835
a2bc16c3
009309df
005300c6
0e560266
00000804
1f540007
101c600c
111c444e
21c34456
179432e4
139c301c
0000311c
60076c0c
301c1294
311c11b4
6c0c0000
12c0101c
0000111c
32e421c3
d0bc0654
009309df
005300c6
08040266
ff96f016
53c340c3
0007c197
600c2a54
444e001c
4456011c
37e470c3
00662294
2254a007
1454c007
139c301c
0000311c
60076c0c
301c1894
311c11b4
6c0c0000
12c0001c
0000011c
37e470c3
01060c54
0ab44067
04c3c037
2abc35c3
009309e0
005300c6
01960086
08040f56
fe967016
10540007
501c800c
511c444e
65c34456
089446e4
80378197
a077a1d7
09e092bc
00c60053
0e560296
00000804
0cd21016
201c600c
211c444e
42c34456
049434e4
09e0b4bc
00c60053
08040856
40c33016
11540007
001c600c
011c444e
50c34456
099435e4
03544047
46f20106
bebc04c3
005309e0
0c5600c6
00000804
50c3f016
62c371c3
58540007
56946687
f5242e24
1250201c
0000211c
6025680c
313c680f
62d24004
301cf324
311c1198
8c0c0000
119c301c
0000311c
40066c0c
54e400b3
910c0554
23e44025
2e24fb14
201cf524
211c1250
680c0000
680f7fe5
4004313c
f32462d2
09f0e4bc
265454e4
0454c027
c00703e6
301c2494
311c11b4
6c0c0000
12c0101c
0000111c
32e421c3
201c1754
211c139c
680c0000
680c69d2
f0ef101c
f0f0111c
32e421c3
05c30935
26c317c3
09e248bc
03860093
02660053
08040f56
1f540007
101c600c
111c5445
21c34d55
179432e4
139c301c
0000311c
60076c0c
301c1294
311c11b4
6c0c0000
12c0101c
0000111c
32e421c3
80bc0654
009309e2
00530386
08040266
40c33016
31540007
001c600c
011c5445
20c34d55
299432e4
14542007
139c301c
0000311c
60076c0c
301c2294
311c11b4
6c0c0000
12c0501c
0000511c
30e405c3
201c1654
211c139c
680c0000
680c6ad2
201c0266
211cf0ef
52c3f0f0
083535e4
f6bc04c3
009309e2
00530386
0c560086
00000804
fd967016
12540007
501c800c
511c5445
65c34d55
0a9446e4
803781d7
a077a217
c0b7c257
09e378bc
03860053
0e560396
00000804
600c0cd2
5445101c
4d55111c
32e421c3
9cbc0494
005309e3
08040386
20c31016
1c540007
001c600c
011c5445
10c34d55
149431e4
139c101c
0000111c
6ad2640c
0266640c
f0ef401c
f0f0411c
31e414c3
02c30635
09e476bc
03860053
08040856
0336f016
50c3ff96
62c381c3
9f5c73c3
00070104
62576254
5f946787
f5242e24
1250201c
0000211c
6025680c
313c680f
62d24004
301cf324
311c1188
8c0c0000
118c301c
0000311c
40066c0c
54e400b3
918c0554
23e44025
2e24fb14
201cf524
211c1250
680c0000
680f7fe5
4004313c
f32462d2
09f0e4bc
2f5454e4
e0070066
c0073154
c2072c54
393c2ab4
36e4108c
301c2614
311c11b4
6c0c0000
12c0201c
0000211c
31e412c3
201c1c54
211c139c
680c0000
680c69d2
f0ef201c
f0f0211c
31e412c3
9f5c0e35
05c30007
26c318c3
debc37c3
00d309e5
00930126
005300a6
01960266
0f56c076
00000804
1f540007
101c600c
111c4555
21c35155
179432e4
139c301c
0000311c
60076c0c
301c1294
311c11b4
6c0c0000
12c0101c
0000111c
32e421c3
1cbc0654
009309e6
00530126
08040266
600c0cd2
4555101c
5155111c
32e421c3
76bc0494
005309e6
08040126
40c33016
25540007
001c600c
011c4555
50c35155
1d9435e4
20070066
40071d54
301c1454
311c139c
6c0c0000
13946007
11b4301c
0000311c
001c6c0c
011c12c0
50c30000
075435e4
c6bc04c3
009309e6
00530126
0c560086
00000804
fd967016
12540007
501c800c
511c4555
65c35155
0a9446e4
803781d7
a077a217
c0b7c257
09e77abc
01260053
0e560396
00000804
600c0cd2
4555101c
5155111c
32e421c3
9ebc0494
005309e7
08040126
40c33016
25540007
001c600c
011c4555
50c35155
1d9435e4
20070066
40071d54
301c1454
311c139c
6c0c0000
13946007
11b4301c
0000311c
001c6c0c
011c12c0
50c30000
075435e4
00bc04c3
009309e8
00530126
0c560086
00000804
0cd21016
201c600c
211c4555
42c35155
049434e4
09e90abc
01260053
08040856
40c33016
25540007
001c600c
011c4555
50c35155
1d9435e4
20070066
40071d54
301c1454
311c139c
6c0c0000
13946007
11b4301c
0000311c
001c6c0c
011c12c0
50c30000
075435e4
14bc04c3
009309e9
00530126
0c560086
00000804
0fd23016
401c600c
411c4d41
54c35345
079435e4
26d26446
09e9cabc
005330c3
03c36186
08040c56
50c3f016
72c361c3
53540007
51946407
f5242e24
1250201c
0000211c
6025680c
313c680f
62d24004
301cf324
311c1180
8c0c0000
1184301c
0000311c
40066c0c
54e400b3
90ac0554
23e44025
2e24fb14
201cf524
211c1250
680c0000
680f7fe5
4004313c
f32462d2
09f0e4bc
215454e4
11b4301c
0000311c
101c6c0c
111c12c0
21c30000
175432e4
139c201c
0000211c
69d2680c
101c680c
111cf0ef
21c3f0f0
093532e4
16c305c3
46bc27c3
009309ea
00530186
0f560266
00000804
1f540007
101c600c
111c4d41
21c35345
179432e4
139c301c
0000311c
60076c0c
301c1294
311c11b4
6c0c0000
12c0101c
0000111c
32e421c3
76bc0654
009309ea
00530186
08040266
00071016
600c2154
4d41201c
5345211c
34e442c3
20071994
301c1454
311c139c
6c0c0000
12946007
11b4301c
0000311c
201c6c0c
211c12c0
42c30000
065434e4
09ead0bc
01860093
00860053
08040856
fe967016
10540007
501c800c
511c4d41
65c35345
089446e4
80378197
a077a1d7
09eb1abc
01860053
0e560296
00000804
600c0cd2
4d41101c
5345111c
32e421c3
38bc0494
005309eb
08040186
0cd21016
201c600c
211c4d41
42c35345
049434e4
09eb9abc
01860053
08040856
600c0cd2
4d41101c
5345111c
32e421c3
a4bc0494
005309eb
08040186
3f36f016
60c3f896
92c321b7
a4d7b3c3
8f5ce517
cf5c02a4
df5c02c4
00070304
0008b2dc
331c6657
64dc00b0
2e240008
201cf524
211c1250
680c0000
680f6025
4004313c
f32462d2
11bc301c
0000311c
373c8c0c
1580fff0
11c0301c
0000311c
61f76c0c
02732006
175464e4
52e4506c
708c0514
5ae4a3c3
02e40f14
508c0514
03e432c3
445c0914
20250444
32c341d7
eb1413e4
a0060053
f5242e24
1250201c
0000211c
7fe5680c
313c680f
62d24004
e4bcf324
64e409f0
a0073f54
19c33f54
3c542007
ec6700a6
01e63c35
001f831c
030638b4
35b4c8e4
d31c0206
31b40001
11b4301c
0000311c
201c6c0c
211c12c0
a2c30000
24543ae4
139c201c
0000211c
69d2680c
101c680c
111cf0ef
21c3f0f0
163532e4
e077a037
00478f5c
0067cf5c
613765d7
00a7df5c
219706c3
3bc329c3
09ebdcbc
01c600d3
00660093
02660053
fc760896
08040f56
139c301c
0000311c
42666c0c
0dd26ff2
101c600c
111c5244
21c35448
059432e4
09ec80bc
005320c3
02c341c6
00000804
0cd21016
201c600c
211c5244
42c35448
049434e4
09ecb4bc
01c60053
08040856
fb967016
16540007
501c800c
511c5244
65c35448
0e9446e4
80378257
a077a297
c0b7c2d7
80f78317
a137a357
09eccabc
01c60053
0e560596
00000804
0136f016
1d540007
401c600c
411c5244
84c35448
159438e4
40078066
301c1354
311c139c
6c0c0000
6cf28266
305c8306
63c304a4
06b416e4
09ed0abc
005340c3
04c381c6
0f568076
00000804
0007f016
600c1a54
5244401c
5448411c
37e474c3
80661294
10544007
23e781e6
301c0db4
311c139c
6c0c0000
66f28266
09ed7ebc
005340c3
04c381c6
08040f56
11b4301c
0000311c
69d26c0c
139c301c
0000311c
63f26c0c
09edf6bc
00000804
1e540007
101c600c
111c5244
21c35448
169432e4
11b4301c
0000311c
101c6c0c
111c12c0
21c30000
0c5432e4
139c301c
0000311c
66f26c0c
09ee36bc
01c60093
02660053
00000804
600c0cd2
5244101c
5448111c
32e421c3
72bc0494
005309ee
080401c6
600c0cd2
5244101c
5448111c
32e421c3
04bc0494
005309f0
080401c6
14540007
101c600c
111c5244
21c35448
0c9432e4
139c301c
0000311c
42666c0c
8ebc66f2
20c309f2
41c60053
080402c3
00077016
600c1654
5244401c
5448411c
36e464c3
80660e94
301c4dd2
311c139c
6c0c0000
66f28266
09f2febc
005340c3
04c381c6
08040e56
600c0cd2
5244101c
5448111c
32e421c3
54bc0494
005309f3
080401c6
600c0cd2
494d101c
4154111c
32e421c3
aabc0494
005309f3
080402a6
00077016
600c1d54
494d401c
4154411c
36e464c3
82c61594
13542007
139c301c
0000311c
82666c0c
f0ef501c
f0f0511c
36e465c3
b8bc06b4
40c309f3
82a60053
0e5604c3
00000804
0336f016
50c3fd96
82c371c3
c31793c3
63540007
65876357
2e246094
201cf524
211c1250
680c0000
680f6025
4004313c
f32462d2
12b8301c
0000311c
301c8c0c
311c12bc
6c0c0000
00b34006
055454e4
4025912c
fb1423e4
f5242e24
1250201c
0000211c
7fe5680c
313c680f
62d24004
e4bcf324
54e409f0
02c63054
60076297
c0272f54
02e60454
2a94c007
11b4301c
0000311c
201c6c0c
211c12c0
12c30000
1d5431e4
139c201c
0000211c
69d2680c
201c680c
211cf0ef
12c3f0f0
0f3531e4
40374297
607762d7
05c3c0b7
28c317c3
c8bc39c3
009309f3
005302a6
03960266
0f56c076
00000804
600c0cd2
494d101c
4154111c
32e421c3
04bc0494
005309f4
080402a6
1f540007
101c600c
111c494d
21c34154
179432e4
139c301c
0000311c
60076c0c
301c1294
311c11b4
6c0c0000
12c0101c
0000111c
32e421c3
50bc0654
009309f4
005302a6
08040266
fe967016
10540007
501c800c
511c494d
65c34154
089446e4
80378197
a077a1d7
09f48cbc
02a60053
0e560296
00000804
236c3016
36542007
f524ae24
6007634c
640c2d54
444e201c
4456211c
34e442c3
40062594
64ac434f
8dd2848c
64af7fe5
648f63f2
438c0113
6baf63ac
40e44f8f
448f0294
60e7618c
305c1194
201c0427
211c1250
680c0000
680f6025
4004353c
f32462d2
09f102bc
353c00b3
62d24004
0c56f324
00000804
50c33016
200641c3
b0bc4506
942f0891
f5240e24
444e301c
4456311c
201c740f
211c1194
280c0000
0010313c
301c680f
311c1190
25f20000
b4cfac0f
00f3b4ef
4cec6c0c
a8cfacef
74cf54ef
4004303c
f32462d2
0c560006
00000804
ae24f016
6006f524
201c600f
211c1194
680c0000
680f7fe5
1190101c
0000111c
640f63f2
40cc0133
68ef60ec
640c4ccf
029430e4
201c440f
211c1250
680c0000
680f6025
6006408c
80ac608f
353c60af
60074004
f3241554
f5240273
6b4f6006
325c6026
ab8c0427
60257c0c
c2d27c0f
02c3f324
09f102bc
25c39fe5
701c0113
711c1250
6e240000
4004633c
1250101c
0000111c
e2948007
f5244e24
7fe5640c
323c640f
62d24004
e4bcf324
000609f0
08040f56
52c3f016
ee2463c3
804cf524
63d2610c
438333e3
0024353c
218324c3
21e463d2
40071894
980f1654
0014353c
60078006
60ac4954
408c68d2
610c46f2
610f31a3
081342c3
404c31e3
604f3283
07538006
615780e6
36546007
11b4301c
0000311c
201c8c0c
211cbecc
534f0013
545c33cf
d3ef0407
40ac136f
0010323c
45f260af
938f808f
00f393af
738f608c
53af4fac
8faf8b8f
718f60e6
51cf4026
726f6157
1250201c
0000211c
6025680c
373c680f
62d24004
04c3f324
09f1a4bc
0424445c
373c00b3
62d24004
04c3f324
08040f56
43c3f016
e197c157
f524ae24
602c23d2
46d2640f
33e3610c
3183204c
83d2680f
700f608c
20acc3d2
e3d2380f
7c0f60cc
4004353c
f32462d2
0f560006
00000804
00000804
f5244e24
323c212f
62d24004
0006f324
00000804
3f36f016
40c3fe96
4e2432c3
f524b2c3
0002341c
14546007
68d260ac
66f2608c
410c31e3
610f32a3
704c0093
704f3183
40043b3c
92dc6007
f324000e
604c1cd3
604f31a3
44d2410c
328331e3
f0ac610f
0007108c
000ce2dc
e027b04c
43cc3694
0404605c
0024363c
158312c3
12e463d2
20072194
63ec1f54
363cac0f
65d20014
504c32e3
704f3283
708f6006
634f70af
0427305c
201cb12c
211c1250
680c0000
680f6025
40043b3c
f32462d2
09f102bc
512c1533
40043b3c
f32462d2
52dc4007
04c3000a
14332664
508f4006
301ca5c3
311c1250
4c0c0000
4c0f4025
c00610c3
6e2496c3
3b3cc3c3
62d24004
bcc3f324
706cf524
400667d2
f0ac506f
a3a3704c
478c10c3
a7cc4037
0404815c
0024d83c
25832ac3
68d23dc3
350332c3
0b0d333c
7f527fe5
658c2383
d31cd3c3
10940007
27544007
4c1167ec
0014383c
35e365d2
3283504c
6006704f
315c674f
478c0427
039412e4
00f30006
6baf67ac
01e44f8f
038c0294
7fe570ac
c5f270af
61c3c78f
00f391c3
62d239c3
40062f8f
91c3478f
2017ffe5
b094e007
710c108f
33e366d2
3283504c
f10f704f
40043c3c
6fd206c3
06c3f324
a38c0193
7c0cf524
7c0f6025
f324c2d2
09f102bc
011305c3
1250701c
0000711c
633c6e24
101c4004
111c1250
00070000
4e24e994
640cf524
640f7fe5
323cb12c
62d24004
e4bcf324
015309f0
706ce4d2
706f6025
3b3cb12c
62d24004
a3d2f324
566404c3
02960006
0f56fc76
00000804
09ecf8bc
09f574bc
00000804
60c3f016
f5242e24
4046e18c
201c418f
211c1250
680c0000
680f6025
4004313c
f32462d2
119c301c
0000311c
301cac0c
311c1198
8c0c0000
704c0213
706c6cd2
099436e4
76bc04c3
706c09e4
039436e4
79f2704c
bfe5910c
2e24b1f2
f98ff524
1250201c
0000211c
7fe5680c
313c680f
62d24004
0f56f324
00000804
436c3016
36544007
f5248e24
6007634c
680c2d54
5445101c
4d55111c
35e451c3
20062594
68ec234f
68ef7fe5
68cf63f2
238c0133
67af63ac
68cc2f8f
029430e4
618c28cf
129461a7
205c43a6
201c0427
211c1250
680c0000
680f6025
4004343c
f32462d2
09f102bc
343c00b3
62d24004
0c56f324
00000804
60c37016
52c341c3
46862006
0891b0bc
b88f982f
f5240e24
5445201c
4d55211c
301c580f
311c1254
201c0000
211cc39c
4c0f0013
119c201c
0000211c
313c280c
680f0010
1198301c
0000311c
cc0f25f2
d92fd90f
6c0c00f3
cd2f4d2c
592fc90f
303c790f
62d24004
0006f324
08040e56
ae24f016
4006f524
201c400f
211c119c
680c0000
680f7fe5
1198101c
0000111c
640f63f2
410c0133
692f612c
640c4d0f
029430e4
206c440f
6027608c
20071694
315c1454
7fe50504
0507315c
315c64f2
01730527
618c416c
4d6f698f
0524315c
039430e4
0527215c
406f4006
1250201c
0000211c
6025680c
40cc680f
60cf6006
60ef80ec
4004353c
15546007
0273f324
6006f524
60266b4f
0427325c
7c0cab8c
7c0f6025
f324c2d2
02bc02c3
9fe509f1
011325c3
1250701c
0000711c
633c6e24
101c4004
111c1250
80070000
4e24e294
640cf524
640f7fe5
4004323c
f32462d2
09f0e4bc
0f560006
00000804
61c37016
f5242e24
11b4301c
0000311c
604c8c0c
25946007
404f4026
608c806f
199432e4
17548007
60af716c
0524245c
698c47d2
0d6f098f
416f618f
045c00b3
016f0527
345c018f
60250504
0507345c
414f4406
4004313c
51546007
09f3f324
54e4a06c
60250994
313c604f
60074004
f3244654
c0070893
301c3b54
311cc418
734f0013
40ec136f
0010323c
45f260ef
938f80cf
00f393af
738f60cc
53af4fac
8faf8b8f
518f41a6
71cf6026
201cd26f
211c1250
680c0000
680f6025
4004313c
f32462d2
6027608c
516c0d94
32e4614c
414f0235
756c316c
043531e4
febc05c3
04c309e3
09f1a4bc
0424045c
313c0133
03a64004
f32465d2
005303a6
0e560006
00000804
0136f016
c1d7a197
8e24e217
f52484c3
802c23d2
43d2840f
280f204c
406c63d2
a3d24c0f
740f60cc
80ecc3d2
e3d2980f
3c0f210c
4004383c
f32462d2
80760006
08040f56
00000804
0736f016
ce2450c3
e0ecf524
07b4e027
4004363c
53546007
0a33f324
e04754cc
2b8c0e94
896c656c
39e494c3
34cf0234
4004363c
43546007
0833f324
0b8c42c3
1250301c
0000311c
40254c0c
54cc4c0f
86c314c3
656c4170
a9e493c3
10c30234
4004363c
f32462d2
f52468c3
079442e4
94c394ec
039479e4
0093038c
0b8cf4ec
02e412c3
42c30354
301cfcd3
311c1250
4c0c0000
4c0f5fe5
0b5410e4
47ac678c
6b8f4faf
078f63ac
2f8f67af
34cf23af
4004383c
f32462d2
09f0e4bc
e0760006
08040f56
0136f016
51c340c3
f5240e24
04e7145c
2fd2318c
345cb16f
35e404c4
71ef0334
b1ef0053
4004303c
60546007
0bd3f324
11b8301c
0000311c
d16c0c10
1250201c
0000211c
6045680c
4066680f
6026518f
326f71cf
4004303c
f32462d2
a4bc04c3
6e2409f1
b16ff524
04c4245c
033425e4
005351ef
341cb1ef
62d20400
04c3f324
09f102bc
f524ee24
11b8001c
0000011c
41e4200c
718c2754
24946007
256c516c
07b421e4
1e9448e4
65e4800f
01331b34
32e471ec
31e41734
800f0cb4
123465e4
301c516c
311c11d0
433c0000
01532b9d
11c8201c
0000211c
31236026
31a3280c
373c680f
62d24004
8076f324
08040f56
0336f016
ce2440c3
404cf524
42dc4007
206c0011
11b4301c
0000311c
50c30c0c
0b5415e4
6047658c
363c0854
60074004
001072dc
2093f324
fff0323c
68d2704f
4004363c
e2dc6007
f324000f
70cc1f73
108c6cf2
106f0af2
4004363c
22dc6007
f324000f
1df370c3
62dc2007
915c000e
708c04a4
39946027
0504315c
315c7fe5
64f20507
0527315c
516c0173
698f718c
315c4d6f
34e40524
215c0394
201c0527
211c1250
680c0000
680f6025
4004363c
f32462d2
0524015c
01b320c3
496c294c
300332c3
0b0d333c
7f5233c4
91e42383
91c30235
ce2454f2
301cf524
311c1250
4c0c0000
4c0f5fe5
602770ec
708c1d35
1a946027
1250201c
0000211c
6025680c
363c680f
62d24004
04c3f324
09e39cbc
ce2470c3
301cf524
311c1250
4c0c0000
4c0f5fe5
e0060053
a007b0cc
201c2b94
211c1250
680c0000
680f6025
4004363c
f32462d2
6027708c
44060a94
106c514f
39e4616c
19c30454
09e3febc
f5242e24
1250301c
0000311c
5fe54c0c
704c4c0f
706f62f2
4004313c
f32462d2
09f0e4bc
708c0c53
0000801c
19946027
356c1070
155c30af
26f20504
0527455c
918f916f
355c0113
4d8c0524
896f8d8f
716f518f
0010313c
0507355c
514f4406
704f6026
70ecb06f
70ef7fe5
70cf63f2
778c00d3
57ac70cf
6b8f4faf
174f0006
0427055c
1250201c
0000211c
6025680c
363c680f
62d24004
708cf324
1a946027
6fd270ec
9cbc04c3
70c309e3
f5246e24
43d250cc
114f096c
0400341c
f32462d2
28d218c3
39e4656c
08c30554
febc19c3
05c309e3
09f102bc
363c0113
62d24004
e3c6f324
e0060053
c07607c3
08040f56
236c3016
3d542007
f5248e24
6007634c
640c3454
4555201c
5155211c
35e452c3
40062c94
656c434f
656f7fe5
654f63f2
438c0133
6baf63ac
654c4f8f
029430e4
618c454f
199460a7
333c648c
7fe50b0d
f88c233c
6d206166
0427305c
1250201c
0000211c
6025680c
343c680f
62d24004
02bcf324
00b309f1
4004343c
f32462d2
08040c56
70c3f016
52c361c3
200643c3
b0bc4786
dc2f0891
153cbc4f
6157100c
2310141d
313c9ccf
7180228d
9d0f7cef
5caf9d2f
0e245c6f
301cf524
311c4555
7c0f5155
118c201c
0000211c
313c280c
680f0010
1188301c
0000311c
ec0f25f2
fdaffd8f
6c0c00f3
edaf4dac
5dafe98f
303c7d8f
62d24004
0006f324
08040f56
ae24f016
6006f524
201c600f
211c118c
680c0000
680f7fe5
1188101c
0000111c
640f63f2
418c0133
69af61ac
640c4d8f
029430e4
201c440f
211c1250
680c0000
680f6025
6006414c
816c614f
353c616f
60074004
f3241554
f5240273
6b4f6006
325c6026
ab8c0427
60257c0c
c2d27c0f
02c3f324
09f102bc
25c39fe5
701c0113
711c1250
6e240000
4004633c
1250101c
0000111c
e2948007
f5244e24
7fe5640c
323c640f
62d24004
e4bcf324
000609f0
08040f56
8e24f016
608cf524
13c364f2
02d353c3
608f6006
60af606c
610f60cc
a16c612f
acd215c3
6006214c
616f614f
1250301c
0000311c
40254c0c
343c4c0f
62d24004
a007f324
41c32b54
701c6e24
711c1250
633c0000
80074004
f5241254
734f6006
0427345c
7c0c938c
7c0f6025
f324c2d2
02bc13ac
bfe509f1
ee94a007
f5242e24
1250201c
0000211c
7fe5680c
313c680f
62d24004
e4bcf324
000609f0
08040f56
0136f016
61c350c3
2e2402c3
f52481c3
74ac356c
61546007
2c942007
744c550c
10c314cc
059421e4
130c333c
007354ec
130c333c
750f6980
7fe574ac
748c74af
748f6025
544c150c
600f780c
40276006
00d304b4
21e13981
60855fe5
55cc5cf2
4004383c
f32462d2
7b544007
266405c3
154c0f13
fff0413c
954f83f2
638c0113
638c754f
43ac754f
6b8f4faf
2006956f
f5cc234f
544c83ec
700f780c
402731c3
00d304b4
31e13981
60855fe5
60065cf2
0427305c
1250201c
0000211c
6025680c
383c680f
62d24004
02bcf324
e00709f1
05c34854
08b37664
3c544007
11b4301c
0000311c
301c8c0c
311ccb38
734f0013
d3efb36f
345c6026
25f20407
938f954f
011393af
738f754c
53af4fac
8faf8b8f
313c954f
756f0010
318f20a6
6026d5cc
126f71cf
1250201c
0000211c
6025680c
383c680f
62d24004
04c3f324
09f1a4bc
0424345c
c3d264f2
666405c3
0424045c
383c0133
01664004
f32465d2
00530166
80760006
08040f56
0136f016
c1d7a197
8e24e217
f52484c3
802c23d2
43d2840f
280f208c
40ac63d2
a3d24c0f
740f614c
816cc3d2
e3d2980f
3c0f218c
4004383c
f32462d2
80760006
08040f56
00000804
0736f016
ce2450c3
e16cf524
07b4e027
4004363c
53546007
0a33f324
e047554c
2b8c0e94
896c656c
39e494c3
354f0234
4004363c
43546007
0833f324
0b8c42c3
1250301c
0000311c
40254c0c
554c4c0f
86c314c3
656c4170
a9e493c3
10c30234
4004363c
f32462d2
f52468c3
079442e4
94c3956c
039479e4
0093038c
0b8cf56c
02e412c3
42c30354
301cfcd3
311c1250
4c0c0000
4c0f5fe5
0b5410e4
47ac678c
6b8f4faf
078f63ac
2f8f67af
354f23af
4004383c
f32462d2
09f0e4bc
e0760006
08040f56
0f36f016
12c361c3
92c34e24
0170f524
600738c3
608c2c94
29546007
204ca10c
423c25c3
980f024f
0d352027
38c341c3
f5810073
9fe5f9e1
9cf26085
100c313c
49807f85
31c320ec
029423e4
410f40cc
602560ac
608c60af
608f7fe5
4004393c
600703c3
000d42dc
0653f324
a007a14c
355c3154
60270404
37ec2d94
e40c404c
6006f80f
04b44027
858100d3
5fe599e1
5cf26085
fff0183c
214f23f2
778c00d3
57ac614f
6b8f4faf
e006216f
755cf74f
201c0427
211c1250
680c0000
680f6025
4004393c
f32462d2
02bc05c3
000609f1
608c13d3
5f546007
5d54a007
204c6110
243c4bc3
580f024f
400631c3
05b42027
7bc30173
f961fd01
40857fe5
313c7bf2
7f85100c
20ec9180
42e421c3
80cc0294
201c810f
211c1250
680c0000
680f6025
7fe5680c
d7ec680f
604ca12c
980c15c3
027f413c
400643c3
04b46027
f9010133
9fe5f561
9cf24085
7f856212
40ec2580
13e432c3
20cc0294
814c212f
fff0183c
214f23f2
738c00d3
53ac614f
6b8f4faf
e006216f
745cf34f
201c0427
211c1250
680c0000
680f6025
4004393c
f32462d2
f39304c3
35542007
11b4301c
0000311c
201c8c0c
211ccb38
534f0013
d3ef136f
345c6006
78c30407
814fe5f2
93af938f
614c00f3
4fac738f
8b8f53af
383c8faf
616f0010
518f40a6
71cf6026
201c326f
211c1250
680c0000
680f6025
4004393c
f32462d2
a4bc04c3
045c09f1
00f30424
4004393c
63d20146
0146f324
0f56f076
00000804
f5244e24
323c21cf
62d24004
0006f324
00000804
0336f016
71c350c3
2e2492c3
f52481c3
60ac216c
2c546007
2a942007
60af7fe5
6025608c
c12c608f
26c3804c
323c7c0c
8027027f
04c30d35
007331c3
39e13d81
60851fe5
343c1cf2
7f85100c
74ec4980
21e413c3
54cc0294
55cc552f
4004383c
f32462d2
7f544007
266405c3
154c0f93
35546007
33540007
fff0413c
954f83f2
638c0113
638c754f
43ac754f
6b8f4faf
2006956f
83ec234f
7c0c544c
31c3700f
04b44027
3d8100d3
5fe531e1
5cf26085
305c6006
95cc0427
1250201c
0000211c
6025680c
383c680f
62d24004
02bcf324
800709f1
05c34854
08b34664
600739c3
301c3b54
311c11b4
8c0c0000
cb38301c
0013311c
b36f734f
6006f3ef
0407345c
954f25f2
93af938f
754c00f3
4fac738f
8b8f53af
313c8faf
756f0010
318f20a6
6026d5cc
327171cf
1250201c
0000211c
6025680c
383c680f
62d24004
04c3f324
09f1a4bc
0424345c
c3d264f2
666405c3
0424045c
383c0133
01664004
f32465d2
00530166
c0760006
08040f56
40c37016
f524ce24
6007608c
604c1694
4004263c
071431e4
40070426
f3243054
05b30426
704f6025
42d270ec
6007f324
04c32554
04533664
133c006c
23f2fff0
00d3306f
706f638c
4faf43ac
308f6b8f
634f6006
0427305c
201cb0ec
211c1250
680c0000
680f6025
4004363c
f32462d2
09f102bc
04c3a3d2
00065664
08040e56
436c3016
36544007
f5248e24
6007634c
680c2d54
4d41101c
5345111c
35e451c3
20062594
688c234f
688f7fe5
686f63f2
238c0133
67af63ac
686c2f8f
029430e4
618c286f
129460c7
205c41a6
201c0427
211c1250
680c0000
680f6025
4004343c
f32462d2
09f102bc
343c00b3
62d24004
0c56f324
00000804
60c37016
52c341c3
44062006
0891b0bc
b84f982f
f5240e24
4d41301c
5345311c
201c780f
211c1184
280c0000
0010313c
301c680f
311c1180
25f20000
d8afcc0f
00f3d8cf
4ccc6c0c
c8afcccf
78af58cf
4004303c
f32462d2
0e560006
00000804
ae24f016
6006f524
201c600f
211c1184
680c0000
680f7fe5
1180101c
0000111c
640f63f2
40ac0133
68cf60cc
640c4caf
029430e4
201c440f
211c1250
680c0000
680f6025
6006406c
808c606f
353c608f
60074004
f3241554
f5240273
6b4f6006
325c6026
ab8c0427
60257c0c
c2d27c0f
02c3f324
09f102bc
25c39fe5
701c0113
711c1250
6e240000
4004633c
1250101c
0000111c
e2948007
f5244e24
7fe5640c
323c640f
62d24004
e4bcf324
000609f0
08040f56
51c33016
f5242e24
6bd2604c
604f7fe5
4004313c
600703c3
f3243c54
07330006
3154a007
11b4301c
0000311c
301c8c0c
311cd414
734f0013
408c136f
0010323c
45f2608f
938f806f
00f393af
738f606c
53af4fac
8faf8b8f
718f60c6
71cf6026
201cb26f
211c1250
680c0000
680f6025
4004313c
f32462d2
a4bc04c3
045c09f1
00f30424
4004313c
63d201a6
01a6f324
08040c56
a157f016
8e24c197
23d2f524
e40fe02c
204c43d2
63d2280f
4c0f406c
608ca3d2
c3d2740f
f80fe0ac
4004343c
f32462d2
0f560006
00000804
00000804
0736f016
ce2450c3
e08cf524
07b4e027
4004363c
53546007
0a33f324
e047546c
2b8c0e94
896c656c
39e494c3
346f0234
4004363c
43546007
0833f324
0b8c42c3
1250301c
0000311c
40254c0c
546c4c0f
86c314c3
656c4170
a9e493c3
10c30234
4004363c
f32462d2
f52468c3
079442e4
94c3948c
039479e4
0093038c
0b8cf48c
02e412c3
42c30354
301cfcd3
311c1250
4c0c0000
4c0f5fe5
0b5410e4
47ac678c
6b8f4faf
078f63ac
2f8f67af
346f23af
4004383c
f32462d2
09f0e4bc
e0760006
08040f56
f5244e24
323c20ef
62d24004
0006f324
00000804
40c37016
f524ce24
6ef2608c
6025604c
40ec604f
4004363c
f32462d2
25544007
266404c3
006c0453
fff0133c
306f23f2
638c00d3
43ac706f
6b8f4faf
6006308f
b0ec634f
0427305c
1250201c
0000211c
6025680c
363c680f
62d24004
02bcf324
a3d209f1
566404c3
0e560006
00000804
1f36f016
81c370c3
a3c392c3
82d7a297
bf5cc317
cf5c01a4
05c301c4
24c33de6
0891b0bc
200607c3
00b0201c
0891b0bc
3e311d51
bc6f5e51
343c9caf
7580fff0
dd6f7c8f
04a7675c
9cf19cd1
175c2406
7df104e7
04c7b75c
5d8f4066
e5c8301c
0013311c
fecf7eaf
101c07c3
111cde38
c4bc0013
0e2409f5
101cf524
111c5244
3c0f5448
11c0201c
0000211c
313c280c
680f0010
11bc301c
0000311c
ec0f27f2
0447775c
0467775c
6c0c0193
0464235c
0467735c
0447725c
0467275c
0447375c
1250201c
0000211c
6025680c
63d7680f
24946027
139c301c
0000311c
80066c0c
101c54c3
111cf0ef
21c3f0f0
0b3532e4
11b8301c
0000311c
54c38c0c
b1ec84d2
71ef716c
4004303c
f32462d2
02bc07c3
800709f1
b1ef1654
303c0293
62d24004
2e24f324
201cf524
211c1250
680c0000
680f7fe5
4004313c
f32462d2
09f0e4bc
f8760006
08040f56
8e243016
618cf524
0b546027
09546047
4004343c
60070226
f3242654
04730226
400f4006
11c0201c
0000211c
7fe5680c
101c680f
111c11bc
63f20000
01b3640f
0444205c
0464305c
0467325c
0447235c
30e4640c
440f0294
4004343c
63d203c3
0006f324
08040c56
f5244e24
0567105c
4004323c
f32462d2
08040006
f5246e24
11b4201c
0000211c
341c080c
62d20400
0804f324
0136f016
c1d7a197
8e24e217
f52484c3
814c23d2
43d2840f
280f218c
402c63d2
a4d24c0f
04a4305c
c4d2740f
04c4405c
e3d2980f
3c0f20cc
44d24257
0444305c
8297680f
238c83d2
383c300f
62d24004
0006f324
0f568076
00000804
11cc301c
0000311c
2c0f2406
1258201c
0000211c
2006680c
4104111c
680f31a3
00000804
41c37016
ce2452c3
305cf524
43e404a4
363c0935
03064004
65546007
0306f324
34e40c53
216c1494
11d0301c
0000311c
1a1d333c
0b9430e4
11c8201c
0000211c
31236026
280c33e3
680f3183
04c4205c
405c540f
305c04c7
43e404e4
81ef0334
61ef0053
11cc301c
0000311c
216cac0c
071451e4
4004363c
34546007
0653f324
071454e4
4004363c
2c546007
0553f324
11b8301c
0000311c
30e46c0c
61ec1f94
0a5431e4
11c8201c
0000211c
31236026
31a3280c
301c680f
311c11d0
201c0000
211c11b8
133c0000
280f5a1d
4004363c
f32462d2
09f0e4bc
363c00b3
62d24004
0006f324
08040e56
0336f016
51c340c3
0e2432c3
245cf524
4c0f04a4
2007318c
545c1454
545c04a7
345c04c7
53e404e4
b16f0434
0073b1ef
71ef716f
4004303c
56546007
0a93f324
518f4066
11b8301c
0000311c
f16ccc0c
1250201c
0000211c
6065680c
6026680f
326f71cf
4004303c
f32462d2
a4bc04c3
545c09f1
545c04a7
345c04c7
53e404e4
b16f0434
0073b1ef
71ef716f
02bc04c3
0e2409f1
301cf524
311c1250
4c0c0000
4c0f5fe5
11b8101c
0000111c
42e4440c
718c1554
12946007
696c3170
98e483c3
46e40db4
840f0b94
083475e4
301c516c
311c11d0
433c0000
303c2b9d
62d24004
e4bcf324
000609f0
0f56c076
00000804
301c3016
311c11b4
2c0c0000
f524ae24
1260301c
0000311c
4c0f44ec
450c856c
0d5421e4
11d0301c
0000311c
4b9d233c
11b8301c
0000311c
4c0f450c
11cc301c
0000311c
04e40c0c
201c0c34
211c11d0
301c0000
311c11b8
423c0000
8c0f0a1d
4004353c
f32462d2
11b8301c
0000311c
31e46c0c
f0bc0354
0c5609f5
00000804
40c31016
f5244e24
11b4301c
0000311c
30e46c0c
323c0794
60074004
f3242b54
618c0533
09546027
07546047
4004323c
20546007
03d3f324
718f6406
4004323c
f32462d2
3de6106c
b0bc50ac
04c30891
de38101c
0013111c
09f5c4bc
f5246e24
318f2066
0400341c
65d203c3
0006f324
04060053
08040856
0336f016
f524ee24
6067618c
301c7a94
311c139c
6c0c0000
61c32006
f0ef201c
f0f0211c
34e442c3
301c0b35
311c11b8
2c0c0000
24d261c3
a56cc5ec
4006a5ef
816c418f
11d0301c
0000311c
4a1d233c
4d944007
4b9d033c
012f010f
11c4801c
0000811c
0001901c
400d393c
540c58c3
28c332a3
301c680f
311c11cc
ac0c0000
48e485c3
8c0f3934
11b8201c
0000211c
63f2680c
0613080f
42e44dec
6d6c2d34
0a5423e4
11c8201c
0000211c
300d393c
31a3280c
301c680f
311c11b8
0c0f0000
4004373c
f32462d2
1250301c
0000311c
301c4c0c
311c139c
8c0c0000
a00642a3
34948007
09f5f0bc
061354c3
0d0f692c
612f092f
51c3410f
c5ef2ad2
00f3a006
a24661ac
400664d2
a32641af
4004373c
f32462d2
11b4301c
0000311c
301c4c0c
311c11b8
8c0c0000
28e484c3
301c0f54
311c1250
4c0c0000
139c301c
0000311c
32a36c0c
f0bc63f2
05c309f5
0f56c076
00000804
301c3016
311c11b4
8c0c0000
f5246e24
0564245c
0400341c
f32462d2
04c344d2
26642006
124c722c
301c3664
311c1254
6c0c0000
04c363d2
2e243664
545cf524
60260564
71cf718f
726f6006
1250201c
0000211c
6025680c
313c680f
62d24004
a4d2f324
202604c3
04c35664
09f1a4bc
08040c56
50c33016
f5244e24
11b4301c
0000311c
87f28c0c
4004323c
3b546007
0733f324
139c301c
0000311c
67d26c0c
4004323c
2f546007
05b3f324
12c0001c
0000011c
41e410c3
323c0794
60074004
f3242254
123c0413
a7f24004
200701c3
f3241b54
031305c3
518f4086
11cf0026
0427345c
301cb26f
311c1250
4c0c0000
4c0f4800
f32422d2
a4bc04c3
045c09f1
00530424
0c560266
00000804
0336f016
4e2470c3
07f2f524
4004323c
50546007
09d3f324
001c600c
011c5244
10c35448
075431e4
4004323c
42546007
0813f324
a7f2bc6c
4004323c
3a546007
0713f324
0544475c
4004323c
600785f2
f3243154
62d205f3
15c3f324
60a004c3
633c6252
363c088c
4580100c
301c2810
311cefef
83c3efef
039498e4
005312c3
c02702c3
0053edb4
680c4085
efef001c
efef011c
31e410c3
6e24f854
25e4f524
24e40535
275c0334
341c0547
62d20400
c076f324
08040f56
00000804
00ff001c
00000804
0136f016
301c40c3
311c11b4
ec0c0000
f524ce24
079447e4
1260301c
0000311c
2c0f30ec
2007318c
000b84dc
518f4066
510c116c
501c712c
511c11d0
24e40000
692f1654
353c4d0f
34e40a1d
253c3a94
101c0b9d
111c11c8
440c0000
31544007
30236026
328333e3
0573640f
0b9d153c
30236026
301c23e3
311c11c4
02c30000
01832c0c
101c0c0f
111c11c8
640c0000
238363d2
501c440f
511c11cc
0ef20000
540f4406
11b8301c
0000311c
363c0c0f
60074004
f3246154
5abc0bf3
140f0a77
11b8101c
0000111c
83c3640c
489448e4
11cc301c
0000311c
301c4c0c
311c11d0
033c0000
040f2a1d
11c8301c
0000311c
00070c0c
201c3554
211c1250
680c0000
680f6025
4004363c
f32462d2
f524ce24
1250201c
0000211c
7fe5680c
5abc680f
301c0a77
311c11d0
233c0000
301c0a1d
311c11cc
6c0c0000
41c329ec
101434e4
11b8301c
0000311c
201c4c0f
211c11c8
60260000
33e33023
3083080c
363c680f
62d24004
301cf324
311c11b8
2c0c0000
72e421c3
301c2254
311c1250
4c0c0000
139c301c
0000311c
42a38c0c
15948007
09f5f0bc
025304c3
fff0313c
60270286
00060735
04542067
71af6026
363c0006
64d24004
0053f324
80760006
08040f56
139c301c
0000311c
301c4c0c
311c1250
6c0c0000
600732a3
301c1094
311c11b4
4c0c0000
11b8301c
0000311c
10c30c0c
035421e4
09f5f0bc
00000804
40c37016
65d2632c
1cbc0985
005309f5
ae24626f
301cf524
311c1250
4c0c0000
4c0f5fe5
718c51cc
5f944007
6a546007
600771ac
718f5694
301c316c
311c11d0
233c0000
40071a1d
433c4694
910f1b9d
201c912f
211c11c4
00260000
100d303c
36a3c80c
301c680f
311c11cc
4c0c0000
16e462c3
2c0f4734
11b8201c
0000211c
63f2680c
07d3880f
12e44dec
6d6c3b34
0a5423e4
11c8201c
0000211c
300d303c
36a3c80c
301c680f
311c11b8
8c0f0000
4004353c
f32462d2
1250301c
0000311c
301c4c0c
311c139c
6c0c0000
600732a3
06b33894
8d0f692c
712f892f
0253510f
006651af
01d3118f
0c546027
0a546047
64f271ac
718f71cf
600600b3
c06671af
301cd18f
311c11b4
4c0c0000
4004353c
f32462d2
11b8301c
0000311c
10c30c0c
0f5421e4
1250301c
0000311c
301c4c0c
311c139c
6c0c0000
63f232a3
09f5f0bc
08040e56
40c3f016
11b4301c
0000311c
47e4ec0c
726c0994
7fe767d2
043c0554
d8bc04c0
ce2409f4
47e4f524
301c0794
311c1260
b0ec0000
201cac0f
211c1250
680c0000
680f7fe5
600771cc
000a92dc
11cf0006
510c316c
001c712c
011c11d0
24e40000
692f1654
303c4d0f
34e41a1d
203c4894
001c1b9d
011c11c8
400c0000
3f544007
31236026
328333e3
0733600f
203c4006
60261b9d
23e33123
11c4301c
0000311c
ac0c02c3
0c0f0583
11c8101c
0000111c
63d2640c
440f2383
11cc501c
0000511c
1a940007
340f2406
11b8301c
0000311c
363c0c0f
62d24004
301cf324
311c1250
4c0c0000
139c301c
0000311c
32a36c0c
6e946007
5abc0d73
140f0a77
11b8101c
0000111c
32c3440c
489443e4
11cc301c
0000311c
301c4c0c
311c11d0
433c0000
840f2a1d
11c8301c
0000311c
00070c0c
201c3554
211c1250
680c0000
680f6025
4004363c
f32462d2
f524ce24
1250201c
0000211c
7fe5680c
5abc680f
301c0a77
311c11d0
233c0000
301c0a1d
311c11cc
6c0c0000
15c3a9ec
101431e4
11b8301c
0000311c
201c4c0f
211c11c8
60260000
33e33023
3483880c
363c680f
62d24004
301cf324
311c11b8
ac0c0000
70e405c3
301c0f54
311c1250
4c0c0000
139c301c
0000311c
32a36c0c
f0bc63f2
0f5609f5
00000804
40c33016
1254301c
0000311c
62d26c0c
043c3664
1cbc04c0
6e2409f5
518cf524
07944047
0400341c
3e546007
0793f324
34544027
0564545c
4004133c
17944007
718f6046
71cf6026
301c526f
311c1250
4c0c0000
4c0f4025
f32422d2
04c3a4d2
56642026
a4bc04c3
03d309f1
518f4046
71cf6026
22d2734c
63d2f324
366404c3
f5246e24
31cf2006
0400341c
f32462d2
04c3a9d2
56642026
341c00b3
62d20400
e4bcf324
000609f0
08040c56
f5244e24
123c618c
60874004
301c0d94
311c1250
4c0c0000
4c0f4025
f32422d2
09f102bc
634c00d3
f32422d2
366462d2
00000804
30c33016
f5240e24
880f8cec
2cef2ccf
11b4201c
0000211c
45c3a80c
069434e4
1260301c
0000311c
303c2c0f
62d24004
0006f324
08040c56
301c3016
311c11b4
2c0c0000
f5240e24
1264301c
0000311c
4c0f4006
25542007
6007658c
44ec2294
301c44cf
311c1260
4c0f0000
21e4450c
656c1854
54c385ec
139435e4
11d0101c
0000111c
3b9d213c
11cc301c
0000311c
301c4c0c
311c11b8
413c0000
8c0f2a1d
4004303c
f32462d2
08040c56
40c31016
f5246e24
4067418c
341c07b4
60070400
f3243d54
033c0773
101c4004
111c1250
40870000
40660f94
6346518f
0427345c
534f4006
6025640c
0007640f
f3241154
606601f3
534c718f
345c6346
640c0427
640f6025
f32402d2
04c343d2
345c2664
63470424
04c30694
09f102bc
01f30006
f5242e24
1250201c
0000211c
7fe5680c
313c680f
62d24004
0366f324
08040856
f5246e24
125c201c
0000211c
341c080c
62d20400
0804f324
810c1016
604c88f2
010566d2
09f4d8bc
005304c3
085602e6
00000804
42c31016
f5244e24
63f2610c
806f204f
4004323c
f32462d2
08560006
00000804
70c3f016
52c341c3
200663c3
b0bc4586
9c2f0891
5c4f4157
7c6f6197
dcafbc8f
f5240e24
494d201c
4154211c
201c5c0f
211c12bc
280c0000
0010313c
301c680f
311c12b8
25f20000
fd2fec0f
00f3fd4f
4d4c6c0c
e92fed4f
7d2f5d4f
4004303c
f32462d2
602761d7
073c0594
d8bc0080
000609f4
08040f56
40c37016
f524ce24
301c010c
311c12a8
4c0c0000
221402e4
12ac301c
0000311c
05e4ac0c
301c1b34
311c12b0
2c0c0000
041401e4
625260a0
612000f3
110c233c
625274a0
233c6980
704c0010
05356207
6d007e05
0053704f
0007504f
143c1654
50cc0080
079412e4
31e4600c
20060c94
0133200f
68af70ec
600c4c8f
039431e4
400f08cf
310f2006
4004363c
f32462d2
0e560006
00000804
40c33016
64d2610c
1cbc0105
0e2409f5
6006f524
201c700f
211c12bc
680c0000
680f7fe5
12b8101c
0000111c
640f63f2
512c0133
694f714c
640c4d2f
029434e4
303c440f
62d24004
0006f324
08040c56
f5242e24
1250201c
0000211c
6025680c
313c680f
62d24004
001cf324
011c12c0
02bc0000
080409f1
0136f016
62c340c3
4e2473c3
f52482c3
602c23d2
c3d2640f
380f2006
504ce3d2
510c5c0f
12a8301c
0000311c
25e4ac0c
301c2414
311c12ac
0c0c0000
1d3420e4
12b0301c
0000311c
21e42c0c
68a00414
00f36252
233c6aa0
60a0110c
69806252
0010233c
6207704c
7e050335
c3d24980
780f6026
5c0fe2d2
23d22197
440f506c
63d261d7
2c0f312c
4004383c
f32462d2
80760006
08040f56
8e243016
400cf524
343c47f2
60074004
f3243a54
5fe70713
343c0794
60074004
f3243254
60cc0613
29946007
fff0323c
02354207
621261e6
12b0201c
0000211c
2e80a80c
12ac301c
0000311c
13e46c0c
65a00a14
3583bf86
12a8201c
0000211c
2e80a80c
45f2440c
00af008f
00d3040f
0c8f68ac
408f08af
20cf60af
4004343c
f32462d2
08040c56
8e243016
20ccf524
13542007
02e4408c
640c0694
30e44006
01130a94
68af60ac
640c4c8f
039430e4
440f28cf
40cf4006
4004343c
f32462d2
08040c56
f5242e24
125c301c
0000311c
313c0c0f
62d24004
0804f324
00ff001c
00000804
00ff001c
00000804
00ff001c
00000804
00ff001c
00000804
00ff001c
00000804
00000804
09f616bc
00000804
00000804
00000804
00000804
00000804
00ff001c
00000804
f5240e24
0ab20804
f3240254
00000804
f9963016
01c05f3c
2054101c
0054111c
fe7e153c
1268201c
0000211c
12a8301c
0000311c
301c4c0f
311c12b0
4c0f0000
efd0201c
0013211c
12ac301c
0000311c
2c0f280c
1110301c
0000311c
848c2c0c
1370301c
0000311c
04ac8c0f
1374301c
0000311c
40060c0f
1378301c
0000311c
650c4c0f
00778037
40f740b7
41774137
12c0001c
0000011c
23c315c3
494d301c
4154311c
09ebdcbc
0c560796
00000804
6006408c
fe7f323c
fe7f123c
4000101c
fe7f123c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
fe7f323c
680f6026
0804404f
139c001c
0000011c
2027200c
08040294
f5242e24
f0160006
03167f36
11b4301c
0000311c
e0510c0c
11b0201c
0000211c
201ce810
211c1260
280c0000
20078006
880f0354
8c0f20cf
0000069c
0e2410c3
08042f24
101cf324
111c11b8
040c0000
140403f2
f524ffb3
11b4101c
0000111c
402c040f
402560cc
201c402f
211c1260
e0500000
8056680f
08940007
fe764056
2ab20f56
f3240254
fe760804
0404ff56
125c101c
0000111c
0025040c
301c040f
311c1260
4c0c0000
0b544007
4c0f5fe5
07944007
1264301c
0000311c
0c0f0026
333c640c
333c00f4
001c100c
011c1268
01800000
4007400c
301c0954
311c1380
00260000
78bc0c0f
301c09f4
311c1380
4c0c0000
1b544027
137c101c
0000111c
0025040c
101c040f
111c12b0
040c0000
301c0085
311c12ac
4c0c0000
069402e4
12a8301c
0000311c
040f0c0c
1264301c
0000311c
40074c0c
1abc0354
080409f3
3f36f016
30c3fd96
494d001c
4154011c
31e410c3
000d34dc
40774006
c01cd2c3
c11c137c
601c0000
611c12b0
701c0000
711c12b4
2e240000
4cc3f524
001c700c
011c125c
400c0000
34e442c3
60251b54
600f0cc3
00f4433c
2f5c8037
001c0001
011c1384
400d0000
621234c3
1268401c
0000411c
780f6e00
60076c0c
0026df54
780c1c0f
40b74c0c
3f3c44d2
68cf0080
4006780c
780c4c0f
0040233c
301c580f
311c12ac
8c0c0000
20e404c3
301c0794
311c12a8
4c0c0000
6006580f
313c7c0f
62d24004
2e24f324
5f3cf524
b1c30040
4004a13c
81c391c3
508c0773
039442e4
00f34006
68af70ac
3f3c4c8f
68cf0080
700c40b7
07356207
700f7e05
908fb0cf
01534006
b070504c
700f702c
b0cf64d2
0053908f
313c70cf
62d24004
43d2f324
26640dc3
f5242bc3
35e470cc
40060b94
3ac350cf
f32462d2
d8bc04c3
29c309f4
323cf524
62d24004
18c3f324
8097f524
c4948007
700c4cc3
125c001c
0000011c
42c3400c
035434e4
1c0f0026
141c1c0c
00070400
301c1e94
311c12c0
40660000
80264d8f
201c8dcf
211c1250
680c0000
680f6e00
1380301c
0000311c
22d20c0f
001cf324
011c12c0
a4bc0000
e89309f1
22dc2007
f324fff4
0396e7f3
0f56fc76
00000804
0f36f016
201cfc96
211c0dbc
3fe60000
29cf29af
1110301c
0000311c
0cf06c0c
01006f3c
363c6006
52c3fc7e
0300b23c
733c6e24
a01c4004
a11c0b84
901c0000
20060001
20772037
1150001c
0000011c
31c326c3
09d8febc
75cc55ac
21832097
40b72383
75ac4df2
20373fe6
1150001c
0000011c
3bc313c3
09d8c8bc
558f0053
758cf524
35cc55ac
21832383
e2d240f7
60d7f324
d6546007
03c360d7
08ce0cbc
436440c3
323c28c3
6dd24a1d
0bb4001c
0000011c
558c3664
400d393c
328333e3
f813758f
1ac30116
0e86640c
80563664
0496f733
0f56f076
00000804
000012a8
006930c3
0c0910c3
c0ac203c
213c2c29
2c49812c
412c013c
00000804
00f7fc96
00612f5c
40d7446d
40b74832
00412f5c
40d7444d
40775032
00212f5c
40d7442d
40375832
00012f5c
0496440d
00000804
400930c3
40874432
01290394
000600b3
029440c7
08040cc9
32c3fe96
32641364
0e946087
1b942227
616b4006
025466a7
123c4026
20770016
00210f5c
60c701f3
22270e94
40060c94
66a762ab
40260254
0016123c
0f5c2037
00530001
02960006
00000804
32c3fe96
32641364
11946087
22942227
214b4006
77a531c3
60273364
40260235
0016123c
0f5c2077
02730021
129460c7
10942227
228b4006
321c31c3
3364fdde
02356027
123c4026
20370016
00010f5c
00060053
08040296
1364fd96
40772364
60873264
40261894
131c40b7
21540806
8006313c
7f327fe5
00574006
202710c3
0f5c0494
20c30021
028303c3
1f5c0037
01d30001
86dd161c
fff0213c
30c30057
003a361c
32837fe5
f88c233c
20b712c3
00413f5c
039603c3
00000804
fe963016
52c31364
32645364
403c6037
608700e0
131c1794
37940800
15c304c3
00013f5c
44bc23c3
402609f8
00074077
04c32e94
3f5c15c3
23c30001
09f81ebc
201c0413
211c86dd
32c30000
1d9413e4
15c304c3
44bc40c6
0ed209f8
1110301c
0000311c
6c0c6c0c
692c4c0c
692f6025
40774026
04c30193
40c615c3
09f81ebc
002602d2
00730077
60776006
00212f5c
029602c3
08040c56
fe963016
301c40c3
311c1110
6c0c0000
06892c0c
60776006
01b323c3
6d01642c
34e44785
60570c54
a02553c3
3f5ca037
60770001
35c3a057
f11430e4
00215f5c
029605c3
08040c56
ff961016
09f8eebc
326430c3
301c6037
311c1110
2c0c0000
0c2c640c
323c4017
618003c7
8f494dcb
341c34c3
68d20001
0504315c
00014f5c
366414c3
315c0113
1f5c05a4
01c30001
366412c3
08560196
00000804
ff96f016
1110601c
0000611c
6c0c780c
eebcac2c
30c309f8
60373264
03c7333c
f1cb9580
32c35209
0001341c
780c6bd2
05c4335c
2f5c04c3
12c30001
00273664
53492554
341c32c3
60070001
104c1354
608903d2
301c6fd2
311c1110
6c0c0000
06c4335c
2f5c05c3
12c30001
366427c3
301c01b3
311c1110
6c0c0000
06e4335c
00012f5c
200602c3
01963664
08040f56
133c30c3
612f3c7f
1780303c
6006614f
602f606f
60cf608f
610f60ef
aaaa301c
aaaa311c
6006604f
01c5305c
600641ef
0804630f
40c3f016
51c362c3
703c5264
301c0980
311c1110
6c0c0000
07c36e2c
36642026
1294a227
05e4345c
c087538b
65850794
0627345c
fc40323c
68050353
0627345c
fb00323c
40060293
1394a0c7
05e4345c
c087538b
67050794
0627345c
fb80323c
698500d3
0627345c
fa40323c
236423c3
0624345c
0587245c
345c6d00
245c0647
32e40604
245c0335
07c30647
08040f56
ff961016
201c40c3
211c0bb4
682c0000
60376dac
60070006
301c2d94
311c1110
6c0c0000
6c6c6c4c
02c36ccc
36642017
20540007
404630c3
347f233c
203c612f
414f2000
406f4017
402f4006
408f4017
6e0040cf
618f616f
410f40ef
aaaa301c
aaaa311c
2f5c604f
205c0001
601701c5
0196630f
08040856
40c37016
eebc61c3
20c309f8
41a72264
4bd20c54
1110301c
0000311c
6c0c6c0c
05d9335c
4e1432e4
f524ae24
05c1245c
245c02c3
323c05c9
045c402c
303c05d1
145c81ac
213c05d9
301cc1ac
311c1110
6c0c0000
0d6c6c0c
21e410c3
353c0735
60074004
f3243154
245c05f3
02c302e1
02e9245c
402c323c
02f1045c
81ac303c
02f9145c
c1ac213c
0321045c
045c10c3
303c0329
145c40ac
313c0331
145c81ac
013c0339
2006c1ac
023520e4
78cc2820
4004253c
043531e4
f32447d2
42d200b3
0026f324
00060053
08040e56
20c31016
226401c3
1110301c
0000311c
2c0c6c0c
03c7323c
4e00842c
31c32b8b
6b8e6025
64d2698c
0f2f69ac
098f0053
085609af
00000804
30c31016
333c3264
082c03c7
0e244c00
8a4bf524
602534c3
694c6a4e
696c64d2
00532c4f
296f294f
4004303c
f32462d2
08040856
0136f016
50c3ff96
326431c3
601c6037
611c1118
580c0000
ec2c680c
006c68ac
30c33664
2e546027
740c380c
04c38d09
243c8d29
0d49402c
812c803c
1f5c84cc
01c30001
123c4d69
546cc42c
10c34664
08540027
6cec780c
00014f5c
366404c3
780c0353
146c6cac
40c33664
13948027
2017780c
03c7213c
1d016d0c
04c33664
40170173
32c348d2
000b361c
033c7fe5
0053f88c
01960026
0f568076
00000804
ae243016
401cf524
411c0bb4
702c0000
72cc4ecc
02c36d2c
702c3664
4ecf4006
4004353c
f32462d2
08040c56
301c7016
311c1110
6c0c0000
305c8c0c
101c02a3
111c9889
21c30000
329432e4
0c4963ec
2e540007
05d9345c
2a1430e4
03c7503c
6e80702c
32c34f49
0008341c
20546007
f524ce24
78bc0146
702c08cc
438b0e80
07944027
218f2006
400621af
0133438e
07354027
2f2c618c
323c218f
638efff0
82bc0146
363c08cc
62d24004
0e56f324
00000804
ff967016
600c50c3
40374006
4cb46047
253c08d3
60c6fa80
0286325c
0bb4301c
0000311c
12c30c0c
08e71abc
602705f3
453c2294
0086f680
08cc78bc
04a4345c
08946027
345c6006
008604a7
08cc82bc
008603b3
08cc82bc
0ef0301c
0000311c
301c4c0c
311c0bb4
0c0c0000
f6c0153c
01932664
0a946047
0bb4301c
0000311c
15c30c0c
e6bc4006
363c08e6
40264004
6ad24037
6026f324
00d36037
f524ce24
c6946007
2f5cf6f3
02c30001
0e560196
00000804
305c1016
600703c1
8e241854
301cf524
311c0bb4
4c2c0000
7ff26acc
00a60acf
301c2066
311c0fe4
4d0c0000
08c8d4bc
4004343c
f32462d2
08040856
51c37016
002c62c3
138c101c
0000111c
089216bc
416440c3
12948007
0bb4301c
0000311c
6c2c6c0c
6c2b6c2c
083560a7
e6bc05c3
04d209f9
04c3180f
00260053
08040e56
f296f016
105c60c3
301c03c1
311c1110
6c0c0000
4c2c6c0c
b2dc2007
313c0012
a98003c7
8007940c
001242dc
0201045c
045c10c3
303c0209
145c40ac
313c0211
245c81ac
323c0219
60a7c1ac
001124dc
04c1145c
145c21c3
313c04c9
245c412c
323c04d1
045c81ac
303c04d9
733cc1ac
07c30e00
c4bc3fe6
36c909d9
5fe521c3
3f5c42f7
63370161
01810f5c
145c16cd
21c30541
0549145c
412c313c
0551245c
81ac323c
0559045c
c1ac303c
2e946007
20072317
245c2b94
02c303a1
03a9245c
402c323c
03b1045c
81ac303c
03b9145c
c1ac213c
2f5c42b7
245c0141
629703c5
420b033c
0f5c0277
045c0121
229703cd
440b213c
2f5c4237
245c0101
629703d5
61f77832
00e10f5c
145c0b73
21c303c1
03c9145c
412c313c
03d1245c
81ac323c
03d9045c
c1ac303c
6c803b8c
2f5c6377
245c01a1
033c03c5
01b7420b
00c11f5c
03cd145c
323c4357
6177440b
00a13f5c
03d5345c
18320357
1f5c0137
145c0081
245c03dd
02c303a1
03a9245c
402c323c
03b1045c
81ac303c
03b9145c
c1ac213c
40f712c3
02c34357
01e431c3
1f5c1b35
145c0061
333c03c5
60b7420b
00410f5c
03cd045c
213c20d7
4077440b
00212f5c
03d5245c
783260d7
0f5c6037
045c0001
145c03dd
21c303c1
03c9145c
412c313c
03d1245c
81ac323c
03d9045c
c1ac203c
03e1145c
145c01c3
313c03e9
045c402c
303c03f1
145c81ac
313c03f9
49a0c1ac
03a1045c
045c10c3
303c03a9
145c40ac
313c03b1
045c81ac
303c03b9
6132c1ac
241423e4
0201245c
245c02c3
323c0209
045c402c
303c0211
145c81ac
313c0219
60a7c1ac
045c1394
10c30221
0229045c
40ac303c
0231145c
81ac313c
245c04c3
123c0239
d6bcc1ac
07c30a0c
09da26bc
0f560e96
00000804
20c37016
a00c61c3
fff0353c
6027204c
001c1cb4
011caaaa
30c3aaaa
109413e4
04a4465c
a0478df2
301c0b94
311c0bb4
0c0c0000
24c312c3
08e6e6bc
365c04d3
600704a4
04331194
aaaa301c
aaaa311c
14e443c3
66bc0494
02f30a40
dddd001c
dddd011c
69ec082f
08cc296c
07946087
0220313c
303c696f
00d3fde0
0360313c
303c696f
68cffca0
08040e56
3f36f016
0f5ce196
21c3035d
00062364
20060777
03dd1f5c
06f70737
1110301c
0000311c
00100c0c
f02c48c3
03591f5c
313c2437
3d8003c7
6e24a40c
f52464f7
34c38749
0001341c
36546007
6007646c
644c3394
2c8964d2
2e542007
0524405c
02013f5c
1f3c03c3
60c606c0
07f24664
873786d7
0001d01c
045305f7
0000d01c
002705f7
00471d54
301c1754
311c1110
6c0c0000
0684435c
20260d66
3f3c42a6
466406b0
34c384d7
0400341c
a2dc6007
f324001a
d01c34f3
df5c0000
153c02e7
24b70180
c537c006
40072dc3
401c1494
411c1110
700c0000
05e4335c
1f3c05c3
36640700
05d760c3
071706d2
0a4066bc
273726d7
03592f5c
03c7323c
47493d80
0014323c
38c36dd2
0121335c
467269d2
4f5c43f7
874d01e1
06370026
20060073
631c2637
159400d7
03594f5c
03c7343c
47493d80
0014323c
05b70026
3a546007
43b74672
01c12f5c
6006474d
065365b7
c5b7c3f2
631c05f3
0e9400d6
03590f5c
03c7303c
2f497d80
300621c3
437721a3
01a12f5c
48c34f4d
cc0f700c
6a4c500c
6a4f6025
00d5631c
301c0c94
311c1110
6c0c0000
0624335c
1f5c05c3
36640359
31c324d7
0400341c
c2dc6007
f3240012
2f5c2533
323c0359
7d8003c7
60076c4c
8c891754
14948007
1110301c
0000311c
335c6c0c
07170644
366415c3
30c304d7
0400341c
e2dc6007
f3240010
18c32173
4717640c
fa80923c
03a79f5c
29c32e71
6a00882b
002bb35c
05770006
03591f5c
03c7313c
604c1d80
19546007
40074c89
60061654
401c6777
411c1110
700c0000
0664435c
2f3c19c3
3f3c0740
466407b0
0f5c0477
05770221
0000b01c
60076757
000c22dc
0382a35c
8fef8c4c
21c33689
313c36a9
56c9412c
81ac323c
103c16e9
2337c1ac
00c0c43c
45942087
01813f5c
0006700d
05c3102d
09f8eebc
326430c3
03d91f5c
41ac213c
2f5c42f7
504d0161
683262d7
0f5c62b7
106d0141
3b3c5031
33640360
1f5c6277
310d0121
62376832
01012f5c
1709512d
172910c3
40ac303c
313c3749
576981ac
c1ac023c
f8bc1cc3
355c09f7
03c30141
0149355c
402c033c
0f5c01f7
114d00e1
283221d7
2f5c21b7
075300c1
700d60c6
102d0006
eebc05c3
30c309f8
1f5c3264
213c03d9
417741ac
00a12f5c
6157504d
61376832
00810f5c
5031106d
04a03b3c
60f73364
00611f5c
6832310d
2f5c60b7
512d0041
24970cc3
b0bc4206
355c08cb
03c30141
0149355c
402c033c
0f5c0077
114d0021
28322057
2f5c2037
516d0001
4c0c38c3
60256a2c
4f5c6a2f
86770359
03c7343c
684c5d80
16946007
31c32b49
0008341c
10546007
1110201c
0000211c
335c680c
4f5c0544
04c30321
36642757
326430c3
05176537
101c0af2
111c1110
640c0000
0484335c
36642757
40074557
fff1a4dc
34c38597
045c48c3
40c30121
326434a3
061765d2
b2dc0007
24d7ffe6
341c31c3
62d20400
1f96f324
0f56fc76
00000804
0f36f016
0f5cf396
21c3015d
00062364
02f70337
1110501c
0000511c
4410340c
6c303ac3
01590f5c
303c0237
0bc303c7
cc0c6180
30c30f49
0001341c
1d546007
0524415c
01011f5c
1f3c01c3
622602c0
04f24664
433742d7
40c306f3
0e540027
0b540047
435c740c
0d660684
42a62026
02b03f3c
14334664
301c8006
311c1110
6c0c0000
0584335c
1f3c06c3
40060300
00073664
2f5c1354
323c0159
1bc303c7
4f496580
500612c3
21f712a3
00e11f5c
2ac32f4d
0c0f680c
86d21013
66bc0317
62d70a40
63176337
fa80833c
08c3ed8a
2dec804c
ad2c21b7
00c0943c
22942087
00c13f5c
0006700d
06c3102d
