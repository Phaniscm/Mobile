768c3664
796c64d2
366405c3
08040e56
205c1016
42c30ab9
0ab1205c
205c42a3
42a30ac1
60ec84d2
36646e6c
085604c3
00000804
60c37016
52c341c3
0fc65364
08cc78bc
300c343c
afcf7980
82bc0fc6
0e5608cc
00000804
60c3f016
842951c3
78bc0fc6
e00608cc
300c343c
54097980
32e46fcc
e0260254
82bc0fc6
07c308cc
08040f56
0736f016
a01c50c3
901c0001
911c0fe4
0bd30000
03c3768c
08ce0cbc
0ee670c3
08cc78bc
8a3c768c
68e3700d
238326c3
0ee6568f
08cc82bc
0280373c
3a1d453c
66127029
21c33580
304e323c
341c3743
6dd20001
341c7069
69f20020
6383680c
31c3c80f
364e233c
4c0f5fe5
341c7069
6ff20008
341c7069
6bf20020
78bc0f06
560c08cc
32a338c3
0f06760f
08cc82bc
341c7069
6fd20002
655c708c
0f200584
0160101c
0011111c
5f7227c3
786c69c3
08745abc
02c35029
340c0065
087348bc
702907f2
002503c3
a2bc340c
768c0872
a1946007
0f56e076
00000804
0136f016
804c71c3
0280313c
3a1d643c
0009865c
300c383c
353cb180
6c0c0700
341c3143
65f20001
20267b2c
03333664
313c15c3
3743304e
0001341c
11946007
6026440c
32a33723
35c3640f
364e233c
4c0f4025
03c37829
300c0025
0872a2bc
341c708c
6ad20001
300c383c
123c5180
6026324e
31a33723
0f06680f
08cc78bc
6026520c
33e33723
720f3283
82bc0f06
807608cc
08040f56
41c33016
313ca04c
233c0020
313c300c
7580300c
135c1501
24c304a4
0fe4301c
0000311c
5abc6c8c
043c0874
340c0030
087348bc
043c06f2
340c0010
0872a2bc
08040c56
0336f016
804c60c3
0001901c
0fe4801c
0000811c
726c0693
0cbc03c3
50c308ce
0280303c
3a1d743c
78bc0ee6
728c08cc
341c3543
67d20001
01c33c29
300c0025
0872a2bc
393c526c
33e3500d
128313c3
528c326f
728f3283
82bc0ee6
04c308cc
2cbc17c3
0ed20880
6c4c7a2c
15c306c3
05c33664
2c6c38c3
0873b4bc
6007726c
c076cb94
08040f56
61c37016
2429a04c
47d200ec
05c360cc
00ff201c
01333664
300c313c
80cc7580
235c05c3
466403a3
03c37829
340c0065
0fe4301c
0000311c
d4bc4d0c
0e5608c8
00000804
0136f016
51c340c3
00f0c04c
646ce429
111c2006
21c37fff
023532e4
7469346f
0008341c
16946007
341c7469
60070020
74691194
0040341c
0ee66df2
08cc78bc
786f784c
82bc0ee6
752c08cc
15c304c3
06c33664
2cbc15c3
09f20880
64cc18c3
342906c3
00ff201c
02b33664
300c373c
6e057980
54096c0c
341c3243
6bd20001
301c0116
311c0b84
6c0c0000
009c001c
80563664
78bc0ee6
5a8c08cc
34098026
100d343c
7a8f32a3
82bc0ee6
04c308cc
301c380c
311c0fe4
4d0c0000
08c8d4bc
0f568076
00000804
0136f016
41c360c3
a04c4364
83c36e24
0f06f524
08cc78bc
e026560c
400d473c
328334e3
79cc760f
06c36dcc
366415c3
82bc0f06
0ee608cc
08cc78bc
43a3766c
0ee6966f
08cc82bc
340c07c3
0fe4301c
0000311c
d4bc4d0c
383c08c8
62d24004
8076f324
08040f56
0086604c
00bc2c0c
08040873
0066604c
00bc2c0c
08040873
0736f016
51c360c3
4230e04c
91c32e24
742cf524
801c67d2
60470000
000934dc
552c0cf3
00ff231c
744c3054
341c3243
60070001
323c2a54
173c0280
756c3a1d
23946047
756f6086
54ec744c
341c3243
6ad20001
0280323c
3a1d373c
0169235c
4d8c55af
672c55cf
202606c3
740c3664
0030033c
d0bc3c0c
393c0872
60074004
000832dc
1013f324
756f6046
54ec744c
341c3243
68f20001
033c740c
3c0c0010
0872a2bc
323c0b33
473c0280
758c3a1d
0001341c
18546007
0644365c
61c76f49
71ac0894
0007341c
3a98001c
02546027
78ec154c
540c2dac
0fe4301c
0000311c
c4bc6c8c
843c0874
604602c0
756c742f
25946047
55af4006
393c55cf
62d24004
74ecf324
1ac36505
06c3440c
3a1d173c
8e242664
4106f524
18c3556f
06c365cc
36642026
033c740c
3c0c0030
0872d0bc
4004343c
28546007
04d3f324
556f4046
01160173
0b84301c
0000311c
001c6c0c
36640082
60068056
740c742f
0030033c
b8bc3c0c
740c0872
0030033c
00bc3c0c
740c0873
0010033c
00bc3c0c
393c0873
62d24004
e076f324
08040f56
0736f016
41c370c3
a04cc40c
81c32e24
742cf524
6087340c
063c0c94
b8bc0010
383c0872
60074004
000b72dc
1693f324
0030a63c
48bc0ac3
0dd20873
0010063c
d0bc340c
383c0872
60074004
000a52dc
1453f324
323c518c
60070014
70ac2294
2d356027
607232c3
301c718f
311c0ba0
4c0b0000
341c32c3
65d20008
7530301c
0093714f
55f0101c
114c314f
26c331ec
0fe4301c
0000311c
5abc6c8c
01f30874
602770ac
32c30cb4
718f6092
301c06c3
311c0fe4
2c8c0000
0873b4bc
512f510c
504c708c
508f2383
63f2708c
708f704c
6007708c
063c1f94
340c0010
0872b8bc
6007760c
760c1154
30cc50cc
21e42383
344c0b94
7cec346f
07c36e4c
04f23664
a2bc340c
383c0872
60074004
f3244554
706c0873
0383104c
0001901c
0cbc0fd2
10ef08ce
39c3306c
33e33023
218323c3
508c506f
708f3283
708c0273
0cbc03c3
10ef08ce
393c508c
33e3000d
708f3283
10c3712c
049431e4
6007708c
712cef94
12c350ec
055431e4
340c0ac3
0872a2bc
6c6c7e0c
40063664
463c542f
04c30010
b8bc340c
04c30872
00bc340c
383c0873
62d24004
e076f324
08040f56
40c37016
605ca04c
560c0644
000675ec
175423e4
6c6c720c
704c3664
4c2f4006
60277829
744c0494
07546047
60277809
744c0794
04946027
355c6006
00260165
08040e56
ff96f016
21c350c3
804c2264
ec6c600c
4047cc2c
245c2694
45d20161
0159345c
16356047
06c37dcc
40662026
30c33664
6ed23264
06c37dcc
40662006
30c33664
66d23264
6d2c760c
366405c3
345c0153
23c30159
40374025
00013f5c
015d345c
0f560196
00000804
105c1016
200703d9
432c1d94
0a544027
18944047
311c6346
6c0b2020
088b033c
66060253
2020311c
01c36c0b
ff00341c
8000101c
0000111c
34e441c3
02c30494
00260053
08040856
fd967016
2046804c
0165145c
0141245c
202512c3
2f5c2077
40b70021
00411f5c
0145145c
62c361cc
4006c412
ac8c4037
363c20c6
56640035
345c6006
0396015d
08040e56
fe967016
145c804c
21c30149
40774025
00211f5c
014d145c
245c4006
61cc0165
0149645c
2006c412
ac8c2037
400620c6
617236c3
40065664
015d245c
0e560296
00000804
ff963016
404c1364
0151325c
a02553c3
3f5ca037
325c0001
325c0155
60470161
325c0e94
31e40141
60860a94
0165325c
6c2c604c
620c64f2
36646c4c
0c560196
00000804
804c1016
0644205c
145c2006
145c018d
145c0195
105c019d
20070361
60261f94
019d345c
233c6b49
341c0034
47d2001c
14946007
145c2026
0213018d
602665d2
0195345c
01160173
0b84301c
0000311c
001c6c0c
366400b5
20268056
01a5145c
0fe4401c
0000411c
20260006
d4bc510c
000608c8
510c2046
08c8d4bc
20660006
d4bc510c
085608c8
00000804
40c37016
205ca04c
746c0644
0001341c
c84c63d2
c86c0053
80bc0106
301c0895
311c0db0
4d090000
255c4dd2
61000584
083436e4
6c6c720c
60063664
0026742f
00060053
08040e56
200600a6
0872a2bc
00000804
fe961016
213401e4
40374006
2fc34077
00403f3c
0875a4bc
111c2e86
640c2200
04c38017
040f03a3
4057040c
308332e3
2085640f
24a3640c
42c322e3
840f4383
640c2085
440f2383
08560296
00000804
60c37016
0cc641c3
08cc78bc
2a548007
0030543c
52835f86
0e64065c
0e84265c
35e46120
82a00514
0e67465c
065c02d3
265c0e24
61200e44
051435e4
465c82a0
01730e27
301c0116
311c0b84
6c0c0000
36640da6
80068056
15c304c3
08cb9cbc
01160153
0b84301c
0000311c
0dc66c0c
80563664
82bc0cc6
04c308cc
08040e56
60c37016
06a4505c
311c6006
4c2b4080
0cab2c6b
54ce8ceb
150e34ee
4d2b952e
0dab2d6b
554e8deb
158e356e
4e4b95ae
0e8b2e6b
55ce8eab
160e35ee
4eeb962e
0f6b2f2b
564e6fab
168e366e
600676ae
4140311c
76ee6c0b
311c6906
6c0b4140
6046770e
4140311c
772e6c0b
03d9365c
2d946007
00471b2c
61860c94
2020311c
77ae6c0b
311c6206
6c0b2020
027377ce
11940027
311c6086
6c0b2020
618677ae
2020311c
77ce6c0b
024a301c
2020311c
77ee6c0b
311c6006
6c0b4105
0206355c
311c6086
6c0b4105
0216355c
0080301c
2100311c
2c2b4c0b
8c8b0c6b
0226255c
0236155c
0246055c
0256455c
2ceb4ccb
6d4b0d2b
0266255c
0276155c
0286055c
0296355c
00a4301c
4105311c
76ce6c0c
311c6006
6c0b4108
02a6355c
311c6506
6c0c4110
02c6355c
08040e56
06a4205c
60062aeb
4140311c
2b0b2c0e
2c0e6905
60464b2b
4140311c
08044c0e
0136f016
007060c3
06a4705c
30e31ccb
40063364
4080211c
1ceb682e
336430e3
1d0b686e
336430e3
1d2b68ae
336430e3
1d4b68ee
336430e3
1d6b692e
336430e3
1d8b696e
336430e3
1dab69ae
336430e3
1e4b69ee
336430e3
1e6b6aee
336430e3
1e8b6b2e
336430e3
1eab6b6e
336430e3
7dcb6bae
9e0b1deb
6a4ebe2b
8a8e0a6e
28c3aaae
01c3688c
366418c3
0223275c
0233175c
0243075c
0253475c
0080301c
2100311c
2c2e4c0e
8c8e0c6e
0263275c
0273175c
0283075c
0293475c
2cee4cce
8d4e0d2e
03d9365c
24946007
00471b2c
5fab0994
311c6186
4c0e2020
60855fcb
002701d3
5fab0d94
311c6086
4c0e2020
61055fcb
5feb4c0e
023e321c
275c4c0e
60060203
4105311c
275c4c0e
60850213
275c4c0e
600602a3
4108311c
275c4c0e
640602c3
4110311c
80764c0f
08040f56
311c6c06
4c0c2200
06a4305c
08044c4f
211c4c06
680c2200
305c65f2
6c4c06a4
0804680f
6c0c610c
20c33664
0084303c
62f20306
323c03c3
63d20014
8003051c
0024323c
051c63d2
323c0180
63d20044
0180051c
0204323c
057262d2
00000804
0084313c
301c6dd2
311c4004
43064128
301c4c0f
311c0408
48064130
313c4c0f
67d20104
0408301c
4130311c
4c0f4406
0014313c
10546007
4004301c
4128311c
8003201c
0000211c
301c4c0f
311c0408
42064130
313c4c0f
60070024
301c1654
311c0418
6c0c4130
0002341c
301c68f2
311c4004
201c4128
4c0f0180
0418301c
4130311c
4c0f4026
0044313c
16546007
0418301c
4130311c
341c6c0c
68f20001
4004301c
4128311c
0180201c
301c4c0f
311c0418
40464130
313c4c0f
67d21004
0418301c
4130311c
4c0f4086
0204313c
301c67d2
311c4004
44064128
313c4c0f
68d20404
0480301c
4130311c
41924c0c
313c4c0f
66d20804
0480301c
4130311c
08046c0c
0014303c
301c67d2
311c0404
42064130
303c4c0f
67d21004
0414301c
4130311c
4c0f4086
0024303c
301c67d2
311c0414
40264130
303c4c0f
67d20044
0414301c
4130311c
4c0f4046
0084303c
301c67d2
311c0404
48064130
303c4c0f
67d20104
0404301c
4130311c
4c0f4406
0404303c
301c68d2
311c0480
4c0c4130
4c0f4172
0804303c
301c66d2
311c0480
6c0c4130
00000804
0014313c
10546007
0404301c
4130311c
4c0f4206
4000301c
4128311c
8023201c
0000211c
313c4c0f
67d21004
0414301c
4130311c
4c0f4086
0024313c
301c6ed2
311c0414
40264130
301c4c0f
311c4000
201c4128
4c0f01a0
0044313c
301c6ed2
311c0414
40464130
301c4c0f
311c4000
201c4128
4c0f01a0
0084313c
301c6dd2
311c0404
48064130
301c4c0f
311c4000
43064128
313c4c0f
67d20104
0404301c
4130311c
4c0f4406
0204313c
301c67d2
311c4000
44064128
313c4c0f
68d20404
0480301c
4130311c
41724c0c
313c4c0f
66d20804
0480301c
4130311c
08046c0c
0014303c
301c67d2
311c0448
44064130
303c4c0f
6fd20024
0448301c
4130311c
4c0f4806
311c6006
201c4140
211c4000
4c0f0003
0044303c
301c68d2
311c0448
201c4130
4c0f0100
0084303c
301c6cd2
311c0448
41064130
60064c0f
4140311c
4c0f4026
0104303c
301c6ed2
311c0448
40864130
60064c0f
4140311c
211c4086
4c0f0100
0204303c
301c6cd2
311c0448
40464130
67064c0f
4140311c
4c0f4406
0404303c
301c67d2
311c0448
42064130
08044c0f
0014303c
301c67d2
311c044c
44064130
303c4c0f
6fd20024
311c6086
201c4140
211c4000
4c0f0003
044c301c
4130311c
4c0f4806
0044303c
301c68d2
311c044c
201c4130
4c0f0100
0084303c
60866cd2
4140311c
4c0f4026
044c301c
4130311c
4c0f4106
0104303c
60866ed2
4140311c
211c4086
4c0f0100
044c301c
4130311c
4c0f4086
0204303c
67866cd2
4140311c
4c0f4406
044c301c
4130311c
4c0f4046
0404303c
301c67d2
311c044c
42064130
08044c0f
0014303c
301c69d2
311c0408
40064130
0001211c
303c4c0f
69d20024
0408301c
4130311c
211c4006
4c0f0010
0044303c
301c69d2
311c0408
40064130
1000211c
303c4c0f
69d20084
0408301c
4130311c
211c4006
4c0f0100
0104303c
301c67d2
311c0418
42064130
08044c0f
003c00e3
003c080d
03640b8d
00000804
0336f016
61c380c3
a04c20f0
75ece429
30430409
0001341c
01166bf2
0b84301c
0000311c
001c6c0c
3664009c
74ac8056
74af7fe5
300c373c
14c39580
304e313c
30431809
0001341c
440c6cd2
30236026
328333e3
34c3640f
364e233c
4c0f5fe5
802655ec
343c3809
33e3100d
75ef3283
78bc0f06
560c08cc
343c1809
33e3000d
760f3283
82bc0f06
373c08cc
f580300c
123c27c3
1809324e
000d343c
318333e3
1809680f
0fe4301c
0000311c
b4bc2c6c
27c30873
384e123c
43237809
318334e3
1809680f
650530c3
153c2006
05c33b9d
2cbc16c3
473c0880
00070080
29c31594
05c368cc
201c3829
366400ff
182973ec
6087340c
00650594
087300bc
002502d3
0872a2bc
73ec0253
0f946107
7fac5809
0b9432e4
301c0116
311c0b84
6c0c0000
009c001c
80563664
588d4006
61ec09c3
366408c3
0f56c076
00000804
70c3f016
402661c3
0ec6448d
08cc78bc
341c7869
60070001
58091194
650532c3
3b9d673c
79acfb4f
fe00201c
0001211c
41e632a3
20db323c
b80979af
78bc0ee6
5eac08cc
343c8026
32a3500d
0ee67eaf
08cc82bc
3c0c04c3
0fe4301c
0000311c
d4bc4d0c
788908c8
0ec67ff2
08cc82bc
08040f56
70c3f016
804c61c3
388d2026
78bc0ec6
0ee608cc
08cc78bc
a026522c
353c3809
32a3100d
0ee6722f
08cc82bc
300c05c3
0fe4301c
0000311c
d4bc4d0c
788908c8
426443c3
0ec69df2
08cc82bc
07c37b2c
366414c3
06c37eec
9cbc2e2c
0f5608cb
00000804
0336f016
50c3ff96
01d091c3
848ce00c
c587d049
c5871d54
c42706b4
c5070754
01331c94
1994c727
620c01b3
30cb6cac
05f33664
686c28c3
366414c3
0361055c
375c02d3
6c2c2784
366424c3
62ac0213
14c36f0c
03b33664
301c0116
311c0b84
6c0c0000
36640ca6
00738056
11540007
0361255c
70cb4af2
28c34037
05c3888c
26c32026
00b34664
4026742c
0245235c
6e4c7c6c
193c07c3
36640040
c0760196
08040f56
0bb4301c
0000311c
48ec4dcc
133c03c3
26640f40
00000804
0336f016
41c360c3
873cee24
901c4004
911c0b84
f5240000
78bc0106
b02c08cc
0106aaf2
08cc82bc
4004373c
24546007
0453f324
62f2700c
7fe51004
702c700f
702f6c0c
704f62f2
82bc0106
28c308cc
f32442d2
01d1355c
79cc67f2
06c36ccc
366415c3
0116fb33
680c29c3
00ad001c
80563664
00a6fa33
b8bc2006
c0760872
08040f56
0f36f016
20b7fd96
b3c34077
01849f5c
28c30010
0cc4a25c
17c4305c
5f866065
201c3283
49a00200
92e469c3
62c30235
2ac36364
fc4fe82c
17c4305c
5f866065
79803283
301c7cce
7c2e00c0
536459c3
17c4305c
32836065
47c37580
606f343c
220604c3
08cb9cbc
353c700c
333c601b
700f232b
275c4006
3f5c0286
704d0041
108d0006
0066b45c
00212f5c
39c351ed
2026af20
313c0393
213c0010
4025080c
003c0ac3
073c2a1d
25c33f9d
0200531c
201c0335
23640200
180c313c
4cce7d80
0010313c
1f5c6037
b5200001
e494a007
0296175c
61cc08c3
17c36cac
03963664
0f56f076
00000804
0bb4201c
0000211c
7f856b2c
04356027
325c6026
301c0587
311c0ba4
6c0c0000
001c6c2c
011c0bb4
36640000
00000804
0037fe96
604730c3
30c32054
1d5460c7
60e730c3
30c31a54
40067f85
60274077
3f5c1635
60770001
32c34017
0f946067
301c0116
311c0b84
6c0c0000
366401e6
40068056
00734077
60776046
00212f5c
029602c3
00000804
60c37016
405c51c3
620c0644
00666e4c
36642026
a6f23089
2af21a0c
00a6628c
1a0c0153
628c25d2
200600a6
628c0093
202600a6
0e563664
00000804
40c37016
0361205c
22944007
513c2c32
c04c0074
600ca8d2
490c4dcc
141c03c3
26640008
6c6c704c
0002341c
10546007
0161365c
0c946087
0116abd2
0b84301c
0000311c
001c6c0c
366400b6
0e568056
00000804
3f36f016
60c3fe96
b05c91c3
a3300de4
0ba4805c
0b0d3d3c
133c7fe5
2077f88c
d31c24f2
07940005
fff4293c
0f0c7aec
0253a800
fff4293c
0002d31c
323c0994
5f860030
5aec3283
ac000b0c
523c00b3
3f860030
796c5183
093c6cec
36641b0b
126410c3
31236026
437223c3
0ba0301c
0000311c
20830c0b
12c342f2
0187313c
265ca3c3
a2840704
8c2b3ac3
0003c35c
796c26f2
06c36dac
366419c3
62200cc3
53e475c3
73c30235
682c2ac3
200606c3
3d3c3664
333c0026
7fe50b0d
f88c233c
605744f2
2f546007
31c32200
027f933c
602f08c3
14544007
00c53b3c
7aec604f
80260f0c
145470e4
0100283c
682f6400
0f0c7aec
3ba37c20
8046684f
3bc30133
273c7272
32a3ffc0
644f18c3
f7a08026
200c343c
698028c3
0080533c
72723bc3
03f36037
08c36200
37c3602f
604f3ba3
1ac3fdd3
06c3642c
36642006
7ce427c3
2cc30235
ffe7055c
05d20057
31c32017
007332a3
3ba332c3
8025740f
a205fd20
e894e007
200c343c
08c37e05
684c4180
6000351c
d31c684f
40540005
61464057
2100311c
0887001c
30944007
0361165c
2e542007
305c182c
60070301
620c2954
0669335c
24546027
341c39c3
331c5000
1e945000
133c62ec
213c00c0
301c804b
311c00f0
4c0e2100
45a062ec
fff4393c
23c36980
301c2364
311c00e4
4c0e2100
311c6146
001c2100
0c0e0487
614600f3
2100311c
0087101c
02962c0e
0f56fc76
00000804
ff963016
505c40c3
432c0ba4
09944047
311c6146
20262020
60c52c0e
00f32c0e
05944027
311c6186
4c0e2020
404743d2
742c0494
742f7f85
65f2732c
6c0c718c
00f33664
059460c7
6c0c71ac
36640086
742c516c
48ec6c0c
1b0b033c
30c32664
333c3264
145c0187
6c800704
04c36c6c
40063664
0587245c
6037732c
15946047
311c6386
6c0b2020
2000341c
2f546007
311c6286
6c0b2020
00f8341c
27946f07
345c6026
03730acd
21c32017
1f944027
111c2006
640b2020
0001341c
17546007
211c4306
680b2020
11946007
640e6017
6dd2680b
00011f5c
0acd145c
0ba4301c
0000311c
6c2c6c0c
366404c3
0c560196
00000804
0ba4301c
0000311c
6c0c6c0c
0bb4001c
0000011c
08043664
a32cf016
0bc4605c
0dc4405c
0894a047
0030313c
3783ff86
0c06305c
a02701b3
313c0894
333c0ff0
323c2a0b
017329ac
105ca3f2
705c0c06
37c30c03
0fff341c
69ac323c
0c06305c
26c314c3
01738006
680f640c
705c644b
37a30e04
8025684f
42052105
75f2644b
200c343c
59807e05
705c684c
37a30e04
6000351c
a8d2684f
311c6346
101c2100
2c0e0287
616c0153
36646c6c
311c6346
201c2100
4c0e0a87
08040f56
40c31016
6007632c
60861794
4010311c
23644c0b
4c0e4172
0361105c
17542007
6e2c602c
12c34da9
323c4dc9
341c40ac
6df20800
60c70113
61ac0694
00466c0c
00b33664
6d6c716c
36642026
66d2732c
00c6704c
00bc2c0c
08560873
00000804
1f36f016
50c3fe96
0704905c
e16c0330
403062d0
0764605c
0361105c
2ac32ad2
435c6a0c
85d20be1
64ec1bc3
1e933664
65d2786c
366405c3
586f4006
355c56ec
055c0da3
8b4c0dc4
428d133c
08cb9cbc
c1c32e24
772cf524
0d9460c7
6c4c75ac
366405c3
3c3c08d2
60074004
000d52dc
1a53f324
0ba0301c
0000311c
34c38c0b
000c341c
13546007
215c19c3
32c30233
0001341c
9e2c6cd2
155c05c3
2f3c0dc4
3fc30040
00274664
00533b54
784c0006
36546047
0056383c
0b0d333c
433c7fe5
84f2f88c
200718c3
7d6c2b94
200605c3
84d23664
6cac756c
758c0073
05c36c2c
20c33664
301c2264
311c0edc
0c2c0000
0361355c
4ed26fd2
4ac30dd2
135c720c
28f20669
0283305c
049460a7
710c4bc3
3c3c3664
60074004
f3247f54
301c0fb3
311c0ba0
4c0b0000
00c4323c
002769d2
5e0c0794
39c3586f
0233635c
323c0773
60070024
493c1454
32c90180
341c31c3
6dd20001
055c7e6c
1f3c0dc4
2fc30040
05d23664
586f5e4c
0493d16b
05c39dcc
0dc4155c
00402f3c
46643fc3
46540007
786f7dec
0edc301c
0000311c
455c0c2c
8ed20361
1ac30dd2
235c660c
48f20669
0283305c
049460a7
650c1bc3
29c33664
cd32c96b
00c6744c
d0bc2c0c
7d6c0872
200605c3
383c3664
6027ffc0
831c0fb4
02940005
74acc026
301c8c0c
0c0c0b00
0dc4155c
466426c3
20570193
831c4017
04940006
6c2c75ac
7d2c0053
366405c3
40043c3c
f32469d2
744c00f3
2c0c00c6
0872b8bc
0296fed3
0f56f876
00000804
fc961016
0e2640c3
08cc78bc
0ef4301c
0000311c
40074c2c
101c1d54
111c0edc
642c0000
644c64d2
00534c2f
101c442f
111c0edc
201c0000
211c0ef4
084c0000
680c044f
6c00040c
2006640f
284f282f
0e26280f
08cc82bc
78bc0e46
301c08cc
311c0f08
4c2c0000
1d544007
0f14101c
0000111c
64d2642c
4c2f644c
442f0053
0f14101c
0000111c
0f08201c
0000211c
644f684c
680c040c
640f6c00
082f0006
080f084f
82bc0e46
0da608cc
08cc78bc
0f20301c
0000311c
60f76c2c
35546007
0f2c201c
0000211c
6007682c
684c1a54
00611f5c
40d72c0d
420b023c
0f5c00b7
0c2d0041
213c20d7
4077440b
00212f5c
00d74c4d
00371832
00011f5c
00732c6d
682f60d7
0f2c101c
0000111c
0f20201c
0000211c
044f084c
040c680c
640f6c00
282f2006
280f284f
82bc0da6
704c08cc
2c0c00c6
0872a2bc
08560496
00000804
60c37016
03c352c3
311c6486
8c0c4600
ffff201c
fe7f211c
24c34283
4c0f5872
36a331c3
32546007
311c6506
2c0c4600
0c0c6a85
4046a0a6
301cc9d2
311c801c
48064113
a0864c0e
31c34006
ffff101c
9fff111c
223c3183
6506e9ac
4600311c
30c34c0f
32835ce6
223c4117
6f8619ac
4600311c
301c4c0f
311c80fc
101c4600
2c0f1c00
500c253c
a0070373
201c1054
211c800c
680c4600
680f6772
0100221c
3f06680c
03a33183
01f3080f
80fc301c
4600311c
1c00201c
203c4c0f
301c500c
311c80f8
4c0f4600
577224c3
311c6486
4c0f4600
08040e56
0ba4105c
236421c3
0080301c
2100311c
213c4c0e
6045808c
205c4c0e
32c30da3
64127fc5
0bc4205c
21c32d00
301c2364
311c0086
4c0e2100
808c213c
4c0e6045
4047432c
61860994
2020311c
4c0e4026
4c0e6085
40270233
60860f94
2020311c
61054c0e
201c4c0e
211c024a
680b2020
66723364
205c680e
49d20361
311c6006
4c0b4105
251c2364
011300f3
311c6006
4c0b4105
251c2364
4c0e00f0
00000804
20267016
03f5105c
0ba4105c
0db3205c
fff0523c
200c353c
323c8580
2580200c
632c306f
07946047
0380301c
a020311c
00d3700f
0080601c
a020611c
9e05d00f
a3d23e05
fdb3bfe5
0bc4405c
0da3305c
ffe0133c
7e056412
313cb180
7180200c
0040233c
632ca84f
07946047
03c0301c
a020311c
00b3680f
611cc806
c80fa020
5e05be05
3fe523d2
105cfdd3
31c30da3
233c7fc5
303c200c
71611800
205c632c
60470da3
323c0a94
6412ffe0
24067180
2020111c
01532c2f
ffe0323c
71806412
0242201c
2020211c
605c4c2f
36c30da3
64127fc5
101c7180
111c8002
2c4f0000
205c4106
20260be7
0da3605c
233c6720
303c230c
716117c0
0da3205c
333c6520
7180230c
611cc086
cc2f4105
0da3205c
333c6520
7180230c
8002601c
0000611c
205ccc4f
65200da3
230c333c
8c6f7180
6c2c614c
0e563664
00000804
6047632c
61460894
2020311c
23c36c0b
01132364
311c6006
6c0b2020
241c23c3
45f2c943
0ac9305c
71546007
0ac9105c
600624d2
0acd305c
6047632c
323c5894
60070044
62063e54
4105311c
101c4c0c
111cffff
2183fff1
4c0f5372
00046006
66676025
201cfd94
211c800c
680c4600
0600351c
4206680f
4105211c
101c680c
111cffff
3183fff1
111c2006
31a3000a
6006680f
60250004
fd946167
211c4206
680c4105
ffff101c
fff1111c
72723183
0004680f
311c6146
40862020
04f34c0e
311c61c6
20262020
61462c0e
2020311c
43462c0e
2020211c
341c680b
7df20004
0380301c
2020311c
01d32c0c
311c6106
40262020
60064c0e
2020311c
63054c0e
13c36c0b
616c1364
36646ccc
00000804
40066006
602541a1
fc9413e4
00000804
60061016
85a200b3
602581a1
5cf25fe5
08040856
21c31016
23e730c3
80061535
8c2e8c0e
8c6e8c4e
8cae8c8e
8cee8cce
8d2e8d0e
8d6e8d4e
8dae8d8e
8dee8dce
3c056405
123cfd73
7c0601f4
01002383
31c320c3
093560e7
880e8006
884e882e
4105886e
fef37f05
0074213c
0184313c
40270180
80060635
016f403c
ff535fc5
08040856
50c33016
209241c3
089168bc
0014343c
760065d2
235c4006
0c56fffd
00000804
31c3ff96
60373064
600648d2
00011f5c
602521a1
fb9423e4
08040196
ff961016
12c331c3
60373064
860743c3
9cbc0494
00d308cb
00013f5c
b0bc13c3
01960891
08040856
0f36f016
a1c390c3
32c362c3
80c36092
e5808384
bc0003c4
8c0038c3
b55c01d3
544b0013
353c346b
700e043f
0016b45c
306e504e
81050105
f2741f27
38c34006
3c008c00
a5620093
4045b141
7fe76800
363cfb74
6ad20014
fff0363c
098029c3
35805ac3
5ebc4026
f0760891
08040f56
08cbeabc
00000804
005330c3
40090025
01a05ef2
00000804
40c33016
600601c3
60250073
41a23364
21e431a2
02c30454
007321c3
02c357f2
0c560120
00000804
ff967016
226440c3
00370006
313c0173
a017008f
a0251282
30e4a037
0c200354
3f5c00d3
32e40001
0006f314
0e560196
00000804
0136f016
70c3fe96
52c361c3
40070006
00d32054
1f542007
50e40025
3c221a54
fbf0813c
00278f5c
00213f5c
632741c3
413c03b4
78220200
fbf0833c
00078f5c
00012f5c
02b44327
43e46405
0073e454
00530006
02961fe6
0f568076
00000804
60061016
88094580
602581a1
88093364
08569af2
00000804
ff963016
400641c3
40250053
7ef26102
00b32100
00015f5c
6025a5a1
a037b182
6180baf2
00011f5c
01962d21
08040c56
51c37016
740910c3
15546007
25c30233
007301c3
40250025
85d28008
63d26808
f95443e4
63f26809
00b301c3
04082025
ee940007
08040e56
0136f016
50c3ff96
815c42c3
28c30000
22544007
0010713c
0ebc07c3
03640892
00530037
740856c3
18546007
16548007
0010653c
38e49fe5
6017f694
24e423c3
06c30db4
3f5c17c3
23c30001
08922abc
00070164
05c3e894
00060053
80760196
08040f56
ff961016
00f330c3
00014f5c
00df433c
5fe52025
840849d2
97f28037
200600b3
00df133c
5cf25fe5
08560196
00000804
40c31016
440c02c3
6980600c
442c700f
323c602c
702f348d
08040856
40c33016
13e40026
000605b4
023542e4
0c560026
00000804
40c31016
440c02c3
69a0600c
442c700f
323c602c
702f350d
08040856
41c33016
13c352c3
043527e7
600f6006
23e702f3
313c0835
343cfe00
600f308d
01d36006
31236026
34837fe5
48a04406
253c3223
32a3108d
343c600f
602f108d
08040c56
40c37016
53c362c3
089326bc
602614c3
7fe53523
44063683
32234aa0
024e213c
640f32a3
08040e56
61c3f016
043563e7
26c312c3
48bc7c05
0f560893
00000804
60c3f016
536451c3
10c30006
711ce006
02138000
373c0112
3483208d
007262d2
02b450e4
402502a0
f5944407
21072085
98810454
fdf34006
08040f56
ff963016
311c6986
40c64140
4c0c4c0f
4c0f4072
305c8026
62f204c1
40068406
098612c3
4140011c
000400b3
00040004
600c0004
511ca006
35830008
523c77d2
a0370010
00012f5c
7392600c
25806332
073424e4
a00fa0c6
6072600c
fd53600f
280c313c
0340141d
0c560196
00000804
40c31016
0084301c
4040311c
61cc2c0b
13646eec
720c3664
4240001c
000f011c
40462ecc
0fe4301c
0000311c
5abc6c8c
08560874
00000804
0136f016
636461c3
13c32264
e28c1264
17c7323c
0564205c
043c8d00
545c0800
35c304b3
345c7fe5
245c04b6
52c30473
fffd541c
0476545c
245c2bd2
345c04e3
23e404f3
35c30514
345c6172
245c0476
c00704d3
0008e2dc
316432c3
04156007
b2dcc047
545c0008
353c0473
60070014
35c31c54
345c6092
145c0476
31c30463
345c6025
345c0466
233c0483
345c0037
32e40433
245c0374
345c0486
345c0483
345c0496
19f304b6
04c6345c
04a3645c
602536c3
236423c3
04a6245c
0413345c
f5dc32e4
245c000b
20070463
145c3754
02c30503
041421e4
0024353c
145c63f2
21e40443
345c1474
23e40443
145c0b74
200704b3
000af4dc
0483245c
04b6245c
323c1533
345c0010
00f30466
0010323c
036403c3
0466045c
8000301c
045c03a3
345c04d6
345c0423
345c0486
345c04b6
a0060496
04a6545c
345c10d3
23e40443
323c0715
23c30010
245c2364
101c0466
21a38000
04d6245c
0423345c
0486345c
04b6345c
0496345c
245c4006
0d7304a6
316432c3
09156007
341c32c3
345c7fff
345c04d6
0bf30466
38542007
0503545c
0463345c
183535e4
0473245c
0024323c
12546007
0466545c
609232c3
0476345c
0423345c
0486345c
04b6345c
0496345c
04a6645c
145c08f3
31c304c3
345c6025
400604c6
04a6245c
0473245c
0014323c
32c369d2
345c6092
60060476
04c6345c
545c0333
35c30493
645c0433
36c304c3
345c6025
145c04c6
245c04a6
323c0473
60070014
32c31054
345c6092
145c0476
345c04c6
345c0423
345c0486
345c04b6
01330496
0493145c
7fe531c3
0496345c
36647c2c
04b3245c
345c45f2
345c0483
807604b6
08040f56
812b3016
2007216b
610b3594
616e612e
604b13c3
0f9413e4
2c948007
65d260cb
60ce7fe5
0313212e
0037213c
32e4606b
03732174
333c40ab
13e40037
323c0554
23c30037
24e42364
60cb1514
7fe569d2
a10b60ce
60eba12e
60ee6072
213c0173
606b0037
067432e4
336432c3
612e610e
0c56616e
00000804
40c33016
00f4203c
170b003c
0fe4301c
0000311c
a0266c2c
323cad21
a006180c
4040511c
68464e80
0047682f
113c0394
280f00a7
00272166
20660554
02940047
80072266
25720215
a00634c3
4000511c
62d23583
282f2272
08040c56
0fe4301c
0000311c
20066c2c
303c2c21
4006180c
4040211c
28466d00
08042c2f
180c303c
211c4006
6d004040
f5244e24
323c0c0c
62d24004
0804f324
301c1016
311c0fe4
8c4c0000
80bc0006
30e30895
0d00504c
08040856
40c31016
0b150007
301c0116
311c0b84
6c0c0000
009e001c
80563664
0fe4201c
0000211c
2c09682c
694c27f2
011c0006
3fe69000
00063664
089580bc
00048220
00040004
00060004
089580bc
60076220
0856f7d4
00000804
101c101c
0000111c
e6bc4386
080408cb
0407105c
408c420f
9ff8101c
ffdf111c
41722183
692c333c
610c608f
0001341c
08047df2
41c31016
101c608c
3183e001
48f2608f
5f26602c
343c3283
602f09ac
20ac01d3
0030323c
080c233c
32236066
318333e3
200d243c
60af32a3
08040856
3f36f016
70c3fd96
42c3a1c3
682c6037
104b833c
d1c32869
000fd41c
28c3a9ab
602c45f2
104bb33c
40ac0133
0030383c
323c6112
b33c308d
712b0034
241c23c3
375c0007
341c0624
68d20008
40676226
5f850635
1100301c
60260053
200dc33c
201c7c8c
3283e000
7c8f6072
233c704c
3b3c084b
7fe50036
f88c933c
42dc4007
2206000c
64f239c3
a83217f3
2ac32106
07c3c82c
38c325c3
d31c6664
09940009
27d219c3
240607c3
38c34006
0895d0bc
ffe03b3c
13b46027
633c708c
cfd225cb
0034563c
a086a2f2
2c303ac3
153c07c3
4006180c
966438c3
fe53daa0
2006706c
0001111c
6cd23183
0624375c
375c7392
2ac30627
07c3684c
28c32066
083c3664
702c680c
0006341c
375c68d2
200604a4
0002111c
00f33183
0484375c
211c4006
32830001
375c67f2
341c0624
60070008
7c8c1254
241c504c
20068000
0028111c
12c342f2
8000201c
07c7211c
351c3283
02330014
504c7c8c
8000241c
111c2006
42f20020
201c12c3
211c8000
328307c7
000c351c
31a330a3
7d0c7c8f
0080341c
702c7df2
0006341c
375c68d2
200604a4
0002111c
00f33183
0484375c
211c4006
32830001
375c66f2
341c0624
64d20008
33647e0c
7e0c00b3
3f5c6077
60b70021
2cc36097
40072383
706c9d94
111c2006
31830001
375c66d2
73720624
0627375c
684c2ac3
1bc307c3
366428c3
101c7c8c
3183e000
7c8f6072
4bd24017
66ac1ac3
366402c3
210600d3
22dc4007
e7d3fff4
03c36097
fc760396
08040f56
0736f016
71c350c3
93c3a2c3
01048f5c
45f228c3
633c602c
0133104b
383c40ac
61120030
308d323c
0034633c
05c39c2c
40c62106
466438c3
684c29c3
0002341c
c0676ad2
9c2c0894
210605c3
00f9201c
466438c3
201c748c
3283e000
748f6072
64d23ac3
0008a31c
9c2c0d94
210605c3
38c34a06
748c4664
e000201c
60723283
e076748f
08040f56
3f36f016
50c3fd96
63c381c3
01c4cf5c
40772364
733c6c2c
5869104b
b41cb2c3
e5f2000f
933c602c
0133104b
373c40ac
61120030
308d323c
0034933c
00c3a65c
60b76006
0615c3e4
7f923cc3
4026c3c3
786c40b7
211c4006
32830001
355c66d2
73720624
0627355c
32c35869
000f341c
28c3e037
05c3888c
23c318c3
466436c3
00863b3c
fff0233c
00363b3c
32a37fe5
f88cd33c
6ed23dc3
882c28c3
210605c3
37c340c6
748c4664
e000201c
60723283
784c748f
084b233c
0036393c
933c7fe5
4007f88c
22065254
65f239c3
aa3c09d3
2106408c
882c28c3
2ac305c3
466437c3
0009b31c
29c30a94
38c348d2
05c38c2c
40062406
466437c3
44f22dc3
60972106
220662d2
341c782c
66d20006
04a4355c
0c4b333c
355c00b3
333c0484
28c30c0b
66d2882c
220605c3
48124057
05c30073
37c34057
748c4664
e000201c
60723283
38c3748f
05c38c6c
26c318c3
46643cc3
4006786c
0001211c
6bd23283
0624355c
355c7392
00b30627
40072106
f613b454
fc760396
08040f56
ff967016
63c350c3
2106842c
46642264
2157748c
241c444c
20068000
0020111c
12c342f2
8000201c
07c7211c
351c3283
363c000c
31a369ac
750c748f
0080341c
b60c7df2
0f5ca037
01960001
08040e56
0336f016
61c340c3
83c392c3
a42ce1d7
40c62106
566437c3
201c708c
3283e000
708f6072
04c3b82c
293c2206
37c3442c
708c5664
e000201c
60723283
c076708f
08040f56
000630c3
1000011c
32e420c3
301c0694
311c0584
00b34130
8584301c
2404311c
001c4c0c
2083ff00
4c0c4c0f
2c0f12a3
00000804
0736f016
71c350c3
400692c3
1000211c
03e432c3
301c0694
311c0584
00b34130
8584301c
2404311c
483c0c10
800700f4
7c4c2694
14c305c3
366429c3
05c39c2c
201c2106
39c300ff
748c4664
e000201c
60723283
7c4c748f
204605c3
366429c3
05c39c2c
201c2106
39c300ff
748c4664
e000201c
60723283
1fd3748f
0804a83c
67d23ac3
707274ac
74ac74af
74af6f72
114b683c
05c37c4c
29c316c3
80273664
000e32dc
16948047
05c39c2c
201c2106
39c300ff
748c4664
e000201c
60723283
9c2c748f
220605c3
ffff201c
0000211c
80670113
9c2c0f94
210605c3
00ff201c
466439c3
201c748c
3283e000
748f6072
80871773
c0070a94
000b72dc
05c39c2c
201c2106
081300f5
0e9480a7
05c39c2c
40c62106
466439c3
201c748c
3283e000
748f6072
80c7fb33
c0071694
0009d2dc
05c39c2c
4cc62106
466439c3
201c748c
3283e000
748f6072
05c39c2c
201c2106
03530099
299480e7
62dcc007
9c2c0008
220605c3
6699201c
466439c3
201c748c
3283e000
748f6072
05c39c2c
201c2206
211c9966
39c30000
748c4664
e000201c
60723283
383c748f
5eac0104
0096001c
064662f2
0c132664
2d948107
211c4006
32c31000
069453e4
311c6346
40064020
301c0173
311c00d4
40064613
301c4c0e
311c00d0
4c0e4613
0104383c
001c5eac
62f20096
26640646
311c6006
23c31000
311c6346
52e44020
301c3354
311c00d4
06134613
30948127
211c4006
32c31000
069453e4
311c6386
40064020
301c0173
311c00e4
40064613
301c4c0e
311c00e0
4c0e4613
0104383c
001c5eac
62f20096
26640646
311c6006
23c31000
00e4301c
4613311c
069452e4
311c6386
42064020
40260053
3ac34c0e
74ac67d2
74af7092
6f9274ac
7c4c74af
200605c3
366429c3
0f56e076
00000804
0136f016
61c350c3
73c382c3
46a661d7
055460a7
61274006
47060254
0002831c
982c1094
210605c3
466437c3
101c748c
3183e000
748f6072
05c3784c
00b318c3
0424365c
16c305c3
366427c3
0f568076
00000804
0f36f016
61c350c3
bf5c72c3
8f5c0124
93c30164
af5c9364
882c0143
210601c3
38c340c6
788c4664
e000201c
60723283
9c2c788f
210606c3
38c329c3
740c4664
111c2006
31830f00
40069c2c
0900211c
31e412c3
06c30494
00732406
210606c3
38c32bc3
9c2c4664
210606c3
38c32ac3
788c4664
e000201c
60723283
740c788f
111c2006
31830f00
211c4006
12c30a00
079431e4
06c39c6c
25c317c3
46646006
0f56f076
00000804
0f36f016
71c360c3
83c392c3
0124bf5c
0144af5c
2106842c
466440c6
201c788c
3283e000
788f6072
06c39c2c
48462106
466438c3
0113a006
06c39c2c
29c32106
466438c3
5be4a025
788cf814
e000201c
60723283
3ac3788f
7eac64d2
36640ac3
0f56f076
00000804
0f36f016
a1c340c3
b3c362c3
833c682c
608c104b
e000101c
60723183
680c608f
a84c2ac3
0034133c
566428c3
933c780c
784c0034
0024233c
4bd2b849
408b333c
220604c3
41ac253c
d0bc38c3
02f30895
ec2c3ac3
0006782c
0007011c
20063083
0001111c
30e401c3
3b3c0594
233c1004
04c3180c
25a32106
766438c3
133c780c
19e4108b
5ac30954
04c3744c
366428c3
933c780c
0ac3108b
582ca02c
200632c3
0007111c
21063183
323c65d2
133c1c0b
04c3180c
38c32bc3
380c5664
341c31c3
60071000
113c1454
19e4120b
5ac30954
04c3744c
366428c3
933c780c
0ac3120b
04c3a02c
40062106
566438c3
2006780c
f000111c
68f23183
4006786c
0780211c
60073283
380c5154
e08c213c
333c786c
733c25cb
113c212c
19e4118b
5ac30954
04c3744c
366428c3
933c780c
780c118b
0800341c
2a946007
67327929
680c283c
3ff4173c
508c073c
708c6cd2
8000501c
07c7511c
a0863583
0028511c
011335a3
501c708c
511c8000
358307c7
32a36272
19ac313c
d9ac303c
710c708f
0080341c
720c7df2
faf2ffe5
573c01f3
a2f20034
0ac3a086
04c36030
180c153c
38c34006
fea0b664
780cf3f2
110b133c
065419e4
744c5ac3
28c304c3
f0763664
08040f56
41c33016
10c353c3
60061364
2100311c
303c2c0e
13c3808c
60462f72
2100311c
14c32c0e
60451364
143c2c0e
6045808c
23642c0e
4c0e6045
201c6085
4c0e8005
a0274106
301c0654
25c30800
4006a3d2
32a36006
0005351c
236423c3
311c6146
4c0e2100
211c41c6
680b2100
0004341c
61c67dd2
2100311c
4c0e4086
08040c56
3f36f016
50c3f896
62c3d1c3
8f5cc3c3
bf5c0264
e5570284
341c602c
61370040
602c6ad2
602f6692
341c750c
7df21000
21372026
341c750c
68f24000
6692742c
750c742f
0400341c
582c7dd2
2004323c
34ac6bf2
104b323c
0040233c
32236026
318333e3
2bc374af
7b8444d2
73833be3
00c78f5c
00e78f5c
980c1b3c
901c20b7
a9c30000
00a79f5c
00103b3c
253c6077
40370400
39c312b3
0001901c
3d946007
2006786c
0001111c
66d23183
0624355c
355c7372
2dc30627
05c3892c
26c31dc3
46643cc3
2006786c
0001111c
60073183
355c1254
73920624
0627355c
133c780c
2177110b
2dc3782c
05c3884c
233c2066
4664104b
101c748c
111c8000
318307c7
557223c3
333c782c
a33c104b
4097692c
780ca2a3
0bcb933c
67327829
805763f2
47c300f3
7ffc731c
401c0335
c4847ffc
42722ac3
3ff4343c
192c233c
508c343c
d92c333c
782c748f
0100341c
001768d2
24c318c3
48bc3bc3
0613089b
0003b31c
24c30e94
341c750c
7df20080
21d7760c
027f313c
5f8521f7
043356f2
0001b31c
24c30e94
341c750c
7df20080
2197760c
016f313c
5fc521b7
023356f2
4ff22bc3
341c750c
7df20080
60f7760c
00613f5c
652118c3
42e44025
8484f494
e007fe20
fff6b4dc
201c748c
3283e000
748f6072
2006786c
0001111c
6ed23183
784c4157
171b323c
782c784f
844c1dc3
12c305c3
104b233c
41174664
602732c3
742c0894
742f6672
341c750c
7dd21000
fc760896
08040f56
341c610c
68f24000
341c608c
7dd20001
6672602c
0804602f
0f36f016
b1c360c3
680c42c3
0400341c
602c64d2
00736472
6492602c
702c782f
011c0006
30830007
111c2006
21c30004
059432e4
0484365c
00937372
0484365c
365c7392
702c0487
0006341c
763c66d2
165c0940
00b304a4
0900763c
0484165c
353cb04c
21c30024
66d25292
78127049
527223c3
106c21a3
8004303c
309212c3
12c363d2
30c33072
2000341c
4d9221c3
21c363d2
30c34d72
1000341c
319212c3
12c363d2
30c33172
4000341c
4e9221c3
21c363d2
30c34e72
8000341c
2f9212c3
12c363d2
706c2f72
25cb333c
08ac133c
0014353c
549221c3
21c363d2
5c0f5472
0080163c
333c702c
333c104b
233c00c7
a1c3100c
363ca284
ed0000c0
323c504c
64d20024
408b323c
70490053
7c0f6812
341c702c
5c0c0200
32c364d2
00736072
609232c3
302c7c0f
44cb313c
10497812
81ac203c
7e32704c
212c233c
333c700c
233c0acb
313c192c
60251c0b
0001341c
092c233c
32a37c0c
500c7c0f
e08c923c
133c704c
702c22cb
08cb833c
0b0b523c
8000241c
8000001c
0002011c
02c342f2
e00c313c
c1ac393c
213c300c
32a3120b
b9ac383c
91ac253c
0034313c
312c233c
108b313c
212c233c
118b313c
112c233c
1ac320a3
706c440f
011c0006
30830001
323c64d2
00f33005
333c700c
333c110b
1ac3412c
b02c640f
341c35c3
331c7000
21547000
1b0b353c
802c0bc3
220606c3
251c23c3
353cc000
4664104b
101c788c
3183e000
788f6072
6572782c
2ac3782f
7c72680c
7c0c680f
011c0006
30a3000c
00937c0f
6592782c
06c3782f
089c92bc
0f56f076
00000804
61c3f016
43c352c3
e1972157
311c6006
59800500
600605f2
0400311c
343c5980
341d0010
03d20130
2c206c80
011387d2
009f423c
00df453c
3bf23fe5
05c304d3
11948027
880b01d3
7c6c800e
411c8006
34830001
402563d2
40450053
00453fc5
027333f2
806705c3
01d31094
800f880c
80067c6c
0001411c
63d23483
00534045
3f854085
33f20085
08040f56
0087f016
00871e54
45c60fb4
8026a006
004765c3
46864c54
49b40047
806640c6
40940027
00c70893
45c61154
8026a686
00c764c3
00e73c14
01070e54
01f33394
a0064746
65c38026
20c30653
8066a686
05b3c026
a7464006
0533c046
81b4301c
4600311c
301c8c0f
311c6000
20064600
60852c0f
60852c0f
60852c0f
60852c0f
60852c0f
60852c0f
60852c0f
60852c0f
60852c0f
60852c0f
321c2c0f
0c0f2198
000606f3
50c320c3
60c38026
111c2006
68802010
080c733c
111c2006
6880104e
100c133c
43644006
016f473c
6472640c
027f313c
40c74025
0087f894
40061935
2010211c
433c7500
2006080c
104e111c
133c7480
4006100c
036406c3
016f043c
6472640c
027f313c
40c74025
0f56f894
00000804
0f36f016
90c3fd96
52c371c3
480c83c3
0304123c
0206313c
b33c7fe5
323cf88c
a01c0034
60670008
361c0754
7fe50002
a33c7f32
7469100c
641c63c3
c0a7000f
c0a73d54
c0470fb4
c0471c54
c00704b4
35f31854
c2dcc067
c0870011
001aa4dc
c10703b3
001152dc
05b4c107
14dcc0e7
1893001a
6654c127
b4dcc147
29f30019
1430740c
20372006
9d0cc077
17c309c3
110b233c
104b383c
2bc30a73
92dc4007
742c0018
104b333c
60373264
09c39cec
47c617c3
0080301c
742c2f73
00370006
9d0cc077
17c309c3
333c4006
4664104b
28f21bc3
4006746c
4000211c
60073283
9c6c1d54
17c309c3
38c325c3
2b3c4664
746c302c
011c0006
30834000
323c68d2
23c3400c
18c34372
81c33f72
00078f5c
09c39cac
35c317c3
540c4664
0034323c
74dc6047
742c0014
20372006
007700a6
09c39d0c
241c17c3
333c0003
4664104b
a01c2713
26070000
744c0694
0bcb333c
0010a33c
0006742c
21260037
9d0c2077
17c309c3
333c4006
4664104b
233c746c
740c25cb
323c7c32
c0c621ac
05356107
6207c046
c0060235
2006746c
4000111c
60073183
9c6c1354
17c309c3
38c325c3
203c4664
38c3400c
60377f72
09c39cac
251c17c3
35c3000f
201c4664
40370300
00266f5c
333c742c
3264104b
9f6c60b7
19c305c3
6e4627c3
60064664
af5c6037
742c0026
104b333c
60b73264
05c39f6c
27c319c3
46646e46
742c1b93
00370006
9d0cc077
17c309c3
333c4006
4664104b
361c744c
333c0400
833c0a8b
740c180c
e08c233c
00c0341c
04946807
100c623c
331c0133
04940080
080c623c
623c0073
742c180c
1b0b233c
333c82a3
3264104b
9cec6037
17c309c3
0081201c
242c363c
cbe64664
2af21bc3
341c740c
601c0030
6207009f
601c0354
742c00df
104b333c
60373264
09c39cec
4c2617c3
742c1213
00370006
9d0cc077
17c309c3
333c4006
4664104b
09c39c6c
25c317c3
466438c3
080c3b3c
41ac203c
00078f5c
09c39cac
35c317c3
540c4664
0034323c
71946047
0006742c
c0770037
09c39d0c
241c17c3
333c0003
4664104b
323c540c
c006e08c
0df46047
311c6006
2383f000
0006c406
3000011c
21e410c3
c6060254
40374006
09c39cec
201c17c3
093300c0
341c744c
801c8000
62f20080
3ac383c3
13546007
0c04323c
623c540c
331ce08c
055400c0
e08c323c
080c633c
0535c107
04b4c207
0053c086
742cc006
00370006
20772146
09c39d0c
400617c3
104b333c
40664664
742c4037
1b0b233c
2b2c223c
00262f5c
104b333c
60b73264
05c39f6c
27c319c3
46646e26
6aa368c3
742cccd2
104b333c
60373264
09c39cec
462617c3
466436c3
341c740c
544c0003
8000241c
42f22086
13a312c3
7b32748c
0444275c
113c09c3
266429ac
f0760396
08040f56
81c0201c
4600211c
6572680c
602c680f
094b333c
201c6812
211c6000
32a311ac
6146640f
7fe50004
201c7ef2
211c81c0
680c4600
680f6592
201c640c
211c6100
328301ac
640c640f
32a34025
0804640f
0736f016
71c350c3
a3c362c3
923c482c
786c104b
144b833c
0006241c
03c68306
0b5440c7
03468206
07544087
01c68106
03544047
01468006
780c342c
134b333c
000d233c
333c782c
233c090b
6066812c
33e33023
23a33183
255c542f
61e60584
33e33423
588c3283
24cb223c
32a32423
0587355c
9c4c782c
200605c3
104b233c
786c4664
211c4006
32830001
0020193c
355c6ad2
63720624
080c213c
200d283c
015332a3
0624255c
080c313c
300d383c
33e36372
355c3283
786c0627
211c4006
32830001
355c66d2
73720624
0627355c
67d23ac3
05c39dcc
26c317c3
46646217
4006786c
0001211c
66d23283
0624355c
355c7392
780c0627
9c4c582c
133c05c3
223c0034
4664104b
4006786c
0800211c
67d23283
06c37fac
27c315c3
00d33664
333c782c
6812094b
786c740f
211c4006
32838000
742c6ad2
742f6772
311c6006
355cfc00
009305a7
6792742c
786c742f
211c4006
32830800
740c64f2
740f6072
23c3748c
782c5972
104b333c
692c333c
786c748f
0200341c
74ac64d2
00736e72
6e9274ac
786c74af
0400341c
74ac64d2
00736f72
6f9274ac
786c74af
0100341c
74ac64d2
00737072
709274ac
782c74af
0c00341c
0400331c
748c0494
00937672
748c64f2
748f7692
4006786c
1000211c
65d23283
0984355c
00936c72
0984355c
355c6c92
7d6c0987
17c305c3
366426c3
341c782c
64d20001
92bc05c3
e076089c
08040f56
0736f016
81c350c3
93c362c3
733c682c
2869104b
441c41c3
602c000f
0040341c
6ad2a3c3
6692602c
750c602f
1000341c
a01c7df2
786c0001
211c4006
32831000
355c66d2
6c920984
0987355c
2006786c
0001111c
66d23183
0624355c
355c7372
28c30627
05c3684c
12c35969
0003141c
366427c3
68d26257
7992748c
750c748f
4000341c
79297df2
6fd26732
06948127
220605c3
06f9201c
05c30093
40c62106
d0bc37c3
02930895
882c28c3
210605c3
37c340c6
784c4664
0002341c
38c369d2
05c38c2c
201c2106
37c300f9
748c4664
e000101c
60723183
784c748f
0002341c
62f22206
931c2106
03940020
00f3596b
00d8931c
590b0394
594b0053
37c305c3
0895d0bc
00c7931c
28c31354
582c882c
200632c3
0007111c
21063183
323c65d2
133c1c0b
05c3180c
37c34217
748c4664
e000201c
60723283
38c3748f
05c38c6c
26c318c3
46646297
2006786c
0001111c
66d23183
0624355c
355c7392
42570627
748c48d2
748f7972
341c750c
7dd24000
0001a31c
742c0894
742f6672
341c750c
7dd21000
2006786c
1000111c
66d23183
0984355c
355c6c72
e0760987
08040f56
3f36f016
50c3f696
72c391c3
02a4df5c
0303cf5c
00b70597
823c482c
3c69104b
341c31c3
61b7000f
c00632c3
0007611c
00063683
0004011c
31e410c3
323c0954
233c1c0b
6026180c
7fe53223
742cd383
0040341c
6ad26137
6692742c
750c742f
1000341c
40267df2
7c6c4137
611cc006
36831000
355c66d2
6c920984
0987355c
00067c6c
0001011c
66d23083
0624355c
355c7372
25970627
bdc32077
af5c21f7
402602e4
600640f7
0c3c6177
0037fff0
29c32573
05c3684c
160b113c
366428c3
67327d29
10546007
63c36197
220605c3
06f9201c
0454c127
210605c3
38c340c6
0895d0bc
09c30293
05c3802c
40c62106
466438c3
341c7c4c
69d20002
842c19c3
210605c3
00f9201c
466438c3
201c748c
3283e000
748f6072
67327d29
11546007
61975d49
05c363c3
c1272106
05c30694
7d892206
41ac223c
d0bc38c3
02530895
982c69c3
210605c3
38c35d49
7c4c4664
0002341c
982c67d2
210605c3
38c35d89
00d74664
23540007
19c37c4c
05c3844c
168b133c
466428c3
882c29c3
32c35c2c
611cc006
36830007
65d22106
1c0b323c
180c133c
2bc305c3
466438c3
30c31d49
00af361c
233c33c4
40f7f88c
c0067c6c
0001611c
6ed23683
0624355c
355c7392
7c4c0627
170b133c
40662177
171b323c
3bc37c4f
3683c017
3ac366f2
0935ace4
00f33cc3
65a01cc3
3ae43364
3ac30235
636463c3
0893c237
09c37c4c
05c3804c
170b133c
466428c3
7c2c54ac
0a4b333c
3e063823
32a32183
465774af
39c34ef2
05c38c2c
61d72106
009f233c
38c361f7
363c4664
0453fff0
10c30657
0e942027
882c29c3
220605c3
233c6057
6077013f
466438c3
ffe0363c
06570233
206710c3
29c30f94
05c3882c
60972406
024f233c
38c360b7
363c4664
63c3ffc0
c0076364
c697bc94
748cc8d2
748f7992
341c750c
7df24000
00067c6c
0001011c
60073083
355c1154
73720624
0627355c
7c4c4157
171b323c
19c37c4f
05c3644c
28c312c3
74ac3664
32835e06
7c0c74af
984c69c3
133c05c3
28c30034
986c4664
19c305c3
38c327c3
06d74664
7aac03d2
26973664
748c28d2
748f7972
341c750c
7dd24000
a2a44217
3c4cb284
c0076ac3
ffed34dc
341c31c3
60078000
01971154
212710c3
05c30694
201c2206
009304fb
210605c3
38c34086
0895d0bc
29c30293
05c3882c
40862106
466438c3
341c7c4c
69d20002
8c2c39c3
210605c3
00fb201c
466438c3
601c748c
3683e000
748f6072
00067c6c
0001011c
66d23083
0624355c
355c7392
21170627
402721c3
742c0894
742f6672
341c750c
7dd21000
c0067c6c
1000611c
66d23683
0984355c
355c6c72
07170987
3c540007
011c0006
10c31000
069451e4
211c4006
42770400
60060173
1200311c
56e463c3
00060594
0800011c
85d70277
01f32006
2dc36257
6c806980
a5976c0c
06c3d481
035430e4
00d30026
9f852085
f1b48067
65970006
01f3ac80
6dc36257
6c807980
32646c09
009f253c
035432e4
00930026
9fe52025
0a9692f2
0f56fc76
00000804
0f36f016
af5cfd96
bf5c0184
8f5c01a4
a82c01c4
0014453c
af5c8af2
bf5c0007
8f5c0027
854c0047
01734664
00078f5c
858c4077
104b053c
2ac313c3
46643bc3
f0760396
08040f56
42c31016
10546007
205c4026
305c0967
341c0964
7cf20001
0624305c
211c4086
32a30004
640c0273
0647305c
233c31c3
205c024e
233c0667
205c024e
6c2c0687
06a7305c
0624305c
305c6272
80070627
700c1154
06c7305c
233c34c3
205c024e
6c2c06e7
0707305c
0624305c
305c6172
08560627
00000804
42c33016
205c53c3
301c0624
31231000
305c32a3
213c0627
323c080c
403c0390
323c3b9d
503c03a0
0c563b9d
00000804
52c33016
610c43c3
0001341c
105c7df2
205c08e7
353c0904
32a3422c
0907305c
6c7260d7
0927305c
08040c56
60c37016
23c342c3
533c6026
0805400d
17544007
07ff231c
790c14b4
0080341c
84d27df2
08948027
60090093
00d3640d
640e600b
600c0073
4aa0640f
fd332680
08040e56
0f36f016
80c3ff96
72c351c3
af5c63c3
63f20144
00d36037
00ff331c
60060a94
9cac6037
17c305c3
38c326c3
0af34664
00f4b33c
801c9bc3
04b30000
05c39c2c
40c62106
46643ac3
201c748c
3283e000
748f6072
05c39c2c
46c62106
46643ac3
05c39c2c
28c32406
46643ac3
201c748c
3283e000
748f6072
311c6006
83840004
ffff921c
400729c3
8b3cda94
c432900c
9c2c0493
210605c3
3ac340c6
748c4664
e000201c
60723283
9c2c748f
210605c3
3ac34726
9c2c4664
240605c3
3ac328c3
748c4664
e000201c
60723283
6006748f
0004311c
dfe58384
dc94c007
f0760196
08040f56
1f36f016
70c3ff96
62c391c3
cf5ca3c3
602c0164
104bb33c
133c606c
400624cb
002682c3
303c00d3
83a3200d
3fe54025
7c0c3bf2
111c2006
31830f00
211c4006
12c30800
189431e4
09c3986c
27c316c3
46643cc3
e03750c3
09c398cc
46a616c3
46643bc3
402c553c
500c283c
538332e3
515c3a3c
400603b3
0a00211c
31e412c3
bf5c0a94
07c30007
26c319c3
3cbc3ac3
02f308a5
09c3986c
27c316c3
46643cc3
100c283c
50c332e3
3a3c5383
53a3115c
0007cf5c
09c398ac
25c316c3
466437c3
f8760196
08040f56
0136f016
50c3fe96
72c361c3
882c83c3
210601c3
60064786
9c2c4664
240606c3
600628c3
740c4664
0003341c
06946047
9c2c742c
220606c3
606700f3
742c0994
06c39c2c
40062406
104b333c
788c4664
041c144c
40068000
0020211c
20c302f2
8000101c
07c7111c
351c3183
32a3000c
790c788f
0080341c
da0c7df2
3f5cc037
60770001
80760296
08040f56
50c3f016
73c361c3
2106842c
46646006
05c3982c
41572106
46646006
341c7c0c
60470003
982c0594
220605c3
606700d3
982c0794
240605c3
32c34006
548c4664
341c7c4c
20068000
0020111c
13c362f2
8000301c
07c7311c
323c2383
31a300c5
750c748f
0080341c
160c7df2
08040f56
0f36f016
50c3fd96
92c3a1c3
608c83c3
608f7672
842c682c
48492106
104b333c
c1064664
b01ce006
750c0006
0080341c
560c7df2
3f5c4077
60b70021
e8d2dfe5
00413f5c
821c28c3
323c0001
c00700df
29c32154
2ac3682c
05c3882c
40062106
104b333c
e0074664
6097e194
5fe523c3
3f5c4037
331c0001
d8b400fd
ef203bc3
00412f5c
821c68c3
263c0001
c02600df
748cf9b3
e000601c
60723683
748c748f
748f7692
039607c3
0f56f076
00000804
30c3ff96
40063264
4010211c
4f85680e
3364680b
00163f5c
00133f5c
0004341c
019678d2
00000804
4f86ff96
4010211c
3364680b
00163f5c
00133f5c
0008341c
600678d2
4010311c
01960c0b
00000804
30c3ff96
40063264
4120211c
4f85680e
3364680b
00163f5c
00133f5c
0004341c
019678d2
00000804
0136f016
50c3ff96
136473c3
436442c3
00e30f5c
01036f5c
11cb313c
70546027
04d46027
71546007
604714f3
60673254
000a34dc
00f4303c
211c4006
61e7f600
60671154
61870354
60260394
361c00b3
7fe50006
233c7f32
0006c00c
f400011c
343c20a3
351c280c
23a3000b
313c540f
69720a4b
200c213c
00ff241c
701232a3
c003351c
343c742f
62520030
0e93744f
00f4303c
211c4006
61e70200
60670d54
61870354
60260394
361c00b3
7fe50006
233c7f32
313cc00c
233c03f4
540fc92c
0104303c
363c67f2
351c280c
23a3000b
05c3540f
211c4006
42a30006
2004313c
722c233c
8004373c
412c133c
027e103c
60076257
31c34154
600f7672
313c07b3
343c00f4
01f329ac
000f141c
343c26f2
351c980c
00f3000a
07942047
900c343c
0014351c
04d3740f
0c942087
200c343c
00a0233c
141d6166
70123230
0037351c
143cfe53
313c180c
416600a0
3320141d
800c033c
06e5303c
341d740f
233c3120
4037fff0
00013f5c
04b46047
806e051c
0006140f
0196142f
0f568076
00000804
63c37016
13640364
11cb303c
28546047
08546067
180c413c
00f4203c
76946027
203c0b93
301c00f4
311cc980
233c0011
313c2d9d
6980180c
141d62a5
303c1320
68d22004
0010313c
0097233c
141d6146
313c1230
6505100c
036403c3
203c0db3
301c00f4
311cc950
233c0011
313c299d
6980180c
141d62a5
403c1320
30c312cb
2000341c
343c68d2
43c3fff0
313c4364
25800014
2004303c
313c68d2
233c0010
61460097
1230141d
100c313c
236423c3
0804303c
343c6df2
62120080
03c36980
66000364
0037333c
780e60c5
343c06b3
62120060
02b36980
c978501c
0011511c
235c6a80
4212ffc1
0160343c
1320341d
2320141d
0010323c
32c322f2
621260a5
036403c3
380e2006
301c02f3
311cc970
ad220011
03944087
200c413c
2004303c
63f24c06
00c0201c
3450141d
03c36980
a0060364
0e56b80e
00000804
ff963016
32c351c3
40063264
001d2f5c
0624105c
07ac40cc
04946027
0524005c
005c0073
3f3c0544
87890040
ffde433c
29858a4c
35c323c3
0f5c4664
01960019
08040c56
ff96f016
20452364
013f613c
0020713c
240b00cc
263c5fe5
4025228d
bc0b4112
830c6037
5d0006c3
466435c3
0f560196
00000804
fe967016
63c340c3
40772264
005ca0cc
145c0624
20070d91
62492754
0014133c
20072037
40571694
62c94432
23e46432
71cc0c94
06056e6c
4b40101c
004c111c
00073664
01131154
00012f5c
009341cd
0002341c
355c69d2
04c30444
00212f5c
26c312c3
02963664
08040e56
0f36f016
72c3ff96
c297a3c3
0624305c
0239935c
009f413c
fff0863c
3e548007
023c4429
640900f4
2d9439e4
208c523c
04d32045
0635c027
8f5c6409
60a70007
af5c0335
a0470007
64090794
b2c34017
0634b3e4
a0270093
64090394
44096037
00013f5c
069423e4
42d76026
e580680f
c02702b3
22250335
22a50053
00071fe5
0153da94
0435c027
0117303c
303c0073
60450157
9fe52580
07c3f853
f0760196
08040f56
ff96f016
72c350c3
0624405c
7a2cc0cc
30c33664
60373064
01c0345c
21c32017
155432e4
00013f5c
01c5345c
255c7269
465c0624
60270484
6b8c0594
2d6c05c3
6b8c0093
2cac05c3
466427c3
0f560196
00000804
205c3016
80cc0624
60276a69
325c1e94
600702a1
313c1a54
60a7fff0
6b8c09b4
912c4bac
0484135c
0444225c
313c0193
60e7ff90
6b8c0ab4
912c4bac
0484135c
0464225c
46646006
08040c56
0f36f016
50c3fe96
01648f5c
936491c3
a364a2c3
60773264
0624705c
7ee9c0cc
60476432
7f8c0754
035c58cc
18c30504
355c2664
6f8c0624
035c58cc
18c30584
8f5c2664
7b700007
19c305c3
4f5c2ac3
34c30021
355cb664
2f8c0624
64327ee9
58cc6705
3a1d013c
266418c3
f0760296
08040f56
fe96f016
207770c3
0544605c
b0cc800c
04c374ac
345c3664
555c0624
04c30444
40062ee9
59ac5664
001c32c3
011cfe00
30830001
35e450c3
7ccc0e54
424b123c
244b223c
00370006
07c38c0c
00215f5c
466435c3
0f560296
00000804
0336f016
21c3fe96
40772264
855ca00c
d4cc0624
0544705c
32c35dac
fe00001c
0001011c
40c33083
345434e4
424b123c
244b223c
00370006
05c33af0
00214f5c
966434c3
00063dac
001e011c
27f21083
0624355c
58cc6f8c
03730fec
211c4006
32c30004
089413e4
0624355c
58cc6f8c
0424035c
800601b3
0002411c
10e404c3
355c0994
6f8c0624
035c58cc
20060404
796c2664
28c305c3
36642969
c0760296
08040f56
1f36f016
c1c3b0c3
07544027
8000901c
2010911c
05944047
8000901c
4103911c
373ce006
1cc3080c
1bc34580
081067a0
233560e7
084c282c
283ca86c
413c808c
603c808c
a53c808c
38c3808c
61123364
4c0e3984
336431c3
39846112
30c38c0e
61123364
cc0e3984
336435c3
39846112
0006a35c
0133e105
808c283c
336438c3
39846112
e0454c0e
cc147be4
0f56f876
00000804
3f36f016
60c3f796
52c341c3
01162bf2
0b84301c
0000311c
001c6c0c
366400d0
c53c8056
35c3e08c
111c2006
31830800
0000a01c
8000a11c
a3c362f2
0cb1265c
1c544007
4007502b
32c31954
241c3164
60077fff
323c0a74
84c3ffc0
ae20201c
0011211c
01938d00
ffc0323c
101c83c3
111cae20
81840011
801c0073
541c0000
a2372000
fff01c3c
2f5c21f7
d2c300e1
3ac3d264
b3c36172
953c54c3
0af3023f
41c3340b
000f441c
46948007
a085f42b
4b54e007
621759cc
31546007
06c3692c
36641ac3
373c59cc
d31c080c
13b40001
bf5c6037
62060027
60f760b7
20666137
81b72177
06c3896c
201c15c3
211c0300
02534103
bf5c6037
62060027
60f760b7
20666137
81b72177
06c3896c
201c15c3
211c1400
60e62010
01534664
06c3692c
36641ac3
15c307c3
50bc2cc3
373c08aa
b580080c
01160153
0b84201c
0000211c
0bc6680c
80563664
ffff921c
600739c3
48c3a894
89c383d2
0996f413
0f56fc76
00000804
30c31016
13c3000b
0ed220c5
fff3315c
401c6212
411c8000
4e004113
ffe3315c
1fe5680e
0856fe53
00000804
ff967016
43c362c3
523c4264
646b0080
2105a037
8cbc4046
163c08cc
800700a0
440b2754
341c32c3
640effcf
31c3396b
03ff341c
34a3940b
fc00241c
740e32a3
41c3392b
001f441c
213c16c3
32c3083e
c000341c
080c033c
343c6f32
980609ac
32a32483
051c640e
18ee1c00
440b0193
351c32c3
640e0030
34c3940b
ff00341c
740e6772
0e560196
00000804
605cf016
5c320624
07544027
8000401c
2010411c
05944047
8000401c
4103411c
0006a46b
6112648b
365c5180
e4ab01c0
33646f80
0045680e
05e42085
0f56f414
00000804
41c33016
343c20cc
60078004
305c1094
a4ec0624
0d91105c
6f8c25d2
0a04135c
6f8c0093
0a24135c
566424c3
08040c56
1f36f016
50c3f696
62c3b1c3
0624805c
65ace0cc
20cb333c
72dc60c7
60c70011
602704b4
13d30b35
d2dc6107
61070026
001bb0dc
f5dc6147
40260030
466d18c3
0104363c
7f4c64f2
366405c3
0024963c
69f239c3
0624355c
9cec6f8c
2dec05c3
466426c3
04c4375c
16c305c3
7dcc3664
1bc305c3
366426c3
0044a63c
80074ac3
355c2394
6f8c0624
0e6c5ccc
259216c3
355c2664
6f8c0624
0c0c5ccc
266416c3
26e918c3
355c2037
4f8c0624
643231c3
323c66a5
4f5c3a1d
28c30001
5ccc8acd
16c303c3
363c2664
6ef20844
0404c75c
1bc305c3
52e948c3
363cc664
64f20084
05c37cac
19c33664
11942007
0624355c
9cec6f8c
2c4c05c3
466426c3
0624355c
9cec6f8c
2c6c05c3
466426c3
40072ac3
355c1d94
6f8c0624
0c2c5ccc
266416c3
6ee938c3
355c60f7
4f8c0624
34c380d7
000f341c
323c6765
2f5c3a1d
18c30061
5ccc46cd
16c303c3
39c32664
34dc6007
355c0028
6f8c0624
0484475c
2d6c05c3
20460e33
326d48c3
0104363c
7f4c63f2
355c3664
6f8c0624
0dec5ccc
266416c3
04c4375c
16c305c3
7dcc3664
1bc305c3
366426c3
0624355c
5ccc6f8c
16c30f2c
26642592
0624355c
5ccc6f8c
16c30f4c
28c32664
41374ae9
0624355c
61174f8c
67056432
3a1d323c
00811f5c
32cd48c3
03c35ccc
266416c3
0624355c
5ccc6f8c
16c30f6c
355c2664
6f8c0624
0fcc5ccc
266416c3
417752e9
0624355c
81574f8c
341c34c3
67c5000f
3a1d323c
00a12f5c
46cd18c3
03c35ccc
266416c3
0624355c
5ccc6f8c
16c30e0c
363c2664
60070024
002124dc
0624355c
475c6f8c
05c30484
26c32cac
40f34664
38c38026
323c8e6d
63f20104
36647f4c
0024a63c
29f21ac3
0624355c
9cec6f8c
2dec05c3
466426c3
04c4375c
16c305c3
7dcc3664
1bc305c3
366426c3
4af22ac3
0624355c
475c6f8c
05c30484
26c32d8c
963c4664
39c30044
23946007
0624355c
5ccc6f8c
16c30e6c
26642592
0624355c
5ccc6f8c
16c30c0c
48c32664
80779309
0624355c
34c34f8c
66a56432
3a1d323c
00212f5c
46cd18c3
03c35ccc
266416c3
0844363c
475c6cf2
05c30404
38c31bc3
36c34f09
375c4664
36640524
8af24ac3
0624355c
9cec6f8c
135c05c3
26c30824
19c34664
355c29f2
6f8c0624
035c5ccc
16c30844
2ac32664
355c4af2
6f8c0624
05c39cec
0864135c
466426c3
69f239c3
0624355c
5ccc6f8c
0884035c
266416c3
930948c3
355c81b7
4f8c0624
341c34c3
6765000f
3a1d323c
00c14f5c
8acd28c3
03c35ccc
266416c3
0624355c
5ccc6f8c
0984035c
266416c3
258918c3
f4dc2007
28c30015
400749a9
0015a2dc
80262a33
8e6d38c3
0104363c
7f4c63f2
a63c3664
1ac30024
355c29f2
6f8c0624
05c39cec
26c32dec
375c4664
05c304c4
366416c3
05c37dcc
26c31bc3
2ac33664
355c4af2
6f8c0624
0484475c
2dac05c3
466426c3
0044963c
600739c3
355c2394
6f8c0624
0e6c5ccc
259216c3
355c2664
6f8c0624
0c0c5ccc
266416c3
930948c3
355c81f7
4f8c0624
643234c3
323c66a5
2f5c3a1d
18c300e1
5ccc46cd
16c303c3
363c2664
6cf20844
0404475c
1bc305c3
4f0938c3
466436c3
0524375c
4ac33664
355c8af2
6f8c0624
05c39cec
0824135c
466426c3
29f219c3
0624355c
5ccc6f8c
0844035c
266416c3
4af22ac3
0624355c
9cec6f8c
135c05c3
26c30904
39c34664
355c69f2
6f8c0624
035c5ccc
16c30924
48c32664
82379309
0624355c
34c34f8c
000f341c
323c6765
4f5c3a1d
28c30101
5ccc8acd
16c303c3
355c2664
6f8c0624
035c5ccc
16c30984
18c32664
20072589
000b04dc
49a928c3
b2dc4007
1453000a
38c38026
363c8e6d
63f20104
36647f4c
0024a63c
29f21ac3
0624355c
9cec6f8c
2dec05c3
466426c3
04c4375c
16c305c3
7dcc3664
1bc305c3
366426c3
4af22ac3
0624355c
475c6f8c
05c30484
26c32dcc
963c4664
39c30044
23946007
0624355c
5ccc6f8c
16c30e6c
26642592
0624355c
5ccc6f8c
16c30c0c
48c32664
80b79329
0624355c
34c34f8c
66a56432
3a1d323c
00412f5c
46cd18c3
03c35ccc
266416c3
0844363c
375c6bf2
05c30444
332948c3
366426c3
0564375c
1ac33664
355c2af2
6f8c0624
05c39cec
0824135c
466426c3
49f229c3
0624355c
5ccc6f8c
0844035c
266416c3
6af23ac3
0624355c
9cec6f8c
135c05c3
26c30944
49c34664
355c89f2
6f8c0624
035c5ccc
16c30964
18c32664
22772729
0624355c
31c34f8c
000f341c
323c6765
2f5c3a1d
18c30121
5ccc46cd
16c303c3
38c32664
6bf26d89
91a948c3
355c88d2
6fac0624
0f0c5ccc
266416c3
f8760a96
08040f56
3f36f016
c0c3bd96
42c32077
00d0d3c3
0624b05c
913c3397
931ce08c
06540001
0002931c
000c94dc
68c30193
0544365c
501c3664
511c8000
101c4103
01530400
305c08c3
36640584
8000501c
4103511c
353c2006
201c6940
4c0e8400
373c75c3
3364023e
3000351c
353c7c0e
c2066420
a53ccc0e
0ac36440
3364600b
402660b7
253c400e
301c6300
680e0080
341c680b
7dd20001
6f3c4006
0f3c08c0
313c00c0
6e80080c
79416c0b
0010313c
6e806112
61416c0b
40452045
0080231c
0006f194
065c6bc3
40060316
0800301c
6f3c2e20
796208c0
033534e4
081431e4
00c00f3c
34e46162
31e40c35
3bc30a34
0313635c
002506c3
3bc30037
0316035c
231c4045
e6940080
64c38006
0f3c24c3
616208c0
03ff331c
321c0335
9180f800
00c01f3c
331c6562
033503ff
f800321c
4045d980
0080231c
931ced94
05940001
315c18c3
00f30524
0002931c
08c30694
0564305c
00b33664
64ac18c3
36640cc3
2ac36097
7c0b680e
cfff341c
253c7c0e
680b2c20
fffe341c
0bc3680e
0313305c
21c32057
18b432e4
f90c343c
003f341c
133c6e00
1de4310c
363c0fd4
341cf90c
6f00003f
2dc46652
067412e4
04d43de4
32e40006
00260d15
28c30173
3664684c
8000501c
2010511c
3000101c
4396e8b3
0f56fc76
00000804
600f6006
00000804
1f36f016
80c3ff96
a2c3b1c3
405ca264
c0cc0624
91c324f2
059371c3
0001a31c
365c0ab4
36640524
0000901c
711ce006
04131000
0003a31c
365c0a94
36640564
0000901c
711ce006
02932000
0448301c
2010311c
18c36c0c
0519115c
202625d2
125c28c3
933c0515
78ac0014
366408c3
51a9e006
e2dc4007
7189000b
a4dc6007
732c000b
732f6025
08958ebc
18c311af
0624215c
0300325c
436443c3
0308525c
8bf2acf2
301c0116
311c0b84
6c0c0000
00c3001c
80563664
0647353c
03156007
00536e20
c3c37180
18c3c164
0624315c
58cc6f8c
04c4035c
266417c3
325c28c3
6fac0624
04c4735c
0080373c
6037bc6b
08c3982c
404613c3
466435c3
60073bc3
a31c1654
04b40001
0544365c
a31c00d3
05940003
0584365c
01333664
0002a31c
19c30694
784c24d2
366408c3
043c9cab
1cbc508b
60c30bfd
32c35ccb
003f341c
200c233c
608c343c
1cbc0980
50c30bfd
1cbc0cc3
20060bfd
42c8111c
0a9584bc
06c330c3
08bc13c3
40c30a95
2cbc14c3
70c30a95
15c305c3
0a952cbc
4000101c
4456111c
0a952cbc
05c360c3
2cbc14c3
101c0a95
111ca000
2cbcc507
30c30a95
13c306c3
0a94a6bc
07c340c3
8000101c
44a4111c
0a952cbc
04c330c3
a6bc13c3
17c30a94
0a9584bc
3bc340c3
a31c68d2
05940002
28c36006
0515325c
10bc2006
04f20a99
411c8006
04c33f80
0a9404bc
00060053
f8760196
08040f56
40c33016
600c51c3
8ebc65f2
100f0895
8ebc0153
20c30895
60a0300c
35e40006
500f0335
0c560026
00000804
0336f016
50c3fe96
91c382c3
605c9264
e0cc0624
e08c323c
04946027
0524375c
604700b3
375c0594
36640564
7cac0073
5b6c3664
6025680c
355c680f
6f8c0624
035c5ccc
18c30664
355c2664
4fac0624
6f8c2a0c
0484335c
0444025c
8f5c0037
9fac0027
402605c3
355c4664
4fac0624
6f8c2a0c
0484335c
0464025c
8f5c0037
9fac0027
404605c3
40264664
02a5265c
08958ebc
19af198f
79ed6006
7472780c
355c780f
2f8c0624
208c393c
5ccc66a5
3a1d013c
266418c3
c0760296
08040f56
3f36f016
60c3ef96
0384cf5c
22f71364
536452c3
62b73264
0624705c
200c20d0
44cc2337
353c4377
7fe50026
53837f52
375c6026
82d702ad
248714c3
24c31054
6c8734c3
b01c0c54
a01cfff8
9f860008
d01c8437
231c0004
09940095
0008b01c
fff8a01c
64376086
fffcd01c
80078297
a0272054
3d3c1e94
6277ffe0
01214f5c
d064d4c3
21c32417
42375fc5
01013f5c
64373064
ffe01a3c
2f5c21f7
a2c300e1
4b3ca064
81b7ffe0
00c11f5c
03f3b1c3
1e94a047
ffd04d3c
1f5c8177
d1c300a1
4417d064
606532c3
4f5c6137
40640081
2a3c8437
40f7ffa0
00613f5c
a064a3c3
00601b3c
2f5c20b7
b2c30041
7ee9b064
63f76432
08958ebc
1daf1d6f
301c0066
311c0fe4
2cac0000
0873b4bc
83b78006
654c2357
36640317
46f24397
4cac7f6c
4caf4025
63970133
802743c3
7f6c0594
40254ccc
365c4ccf
4e6b0624
0143835c
20066e4b
19c32037
0464415c
12c306c3
466428c3
12dc0007
4397000e
602532c3
602763b7
7e290694
d9dc6027
2113000a
32c34397
22946047
4cec7f6c
4cef4025
01c14f5c
23d79e2d
404721c3
365c0a54
6f8c0624
50cc49c3
0524035c
26641cc3
061019c3
a04725c3
40060254
0007cf5c
82d706c3
1d8414c3
239702b3
406721c3
7f6c1694
40254d0c
39c34d0f
25c30e10
0254a047
cf5c4006
06c30007
841762d7
4f5c2e00
34c30141
0db38664
21c32397
1e944087
4d2c7f6c
4d2f4025
62d7acf2
431c43c3
079400c4
0d89165c
439724d2
a5c342f7
0e1039c3
a04725c3
40060254
0007cf5c
62d706c3
1a8413c3
2397fb73
40a721c3
7f6c1e94
40254d4c
acf24d4f
43c362d7
08948107
0d89165c
301c25d2
62f700c8
49c3b5c3
25c31210
0254a047
cf5c4006
06c30007
13c362d7
f7531b84
21c32397
279440c7
696c5f6c
696f6025
7e2d6066
0007cf5c
121049c3
42d706c3
25c312c3
01414f5c
866434c3
0624265c
0229325c
03546027
06946127
24c66006
4020111c
6b8c640e
50cc49c3
0544035c
26641cc3
0624365c
19c36f8c
035c44cc
1cc30584
43972664
60c732c3
fff1a4dc
0624265c
0229325c
03546027
06946127
311c64c6
80864020
6b8c8c0e
44cc19c3
0564035c
26641cc3
8238301c
2010311c
0f0f201c
00f34c0e
43c36397
03b48027
3e2d2026
40043c3c
60076077
4f5c1594
9ead0161
3e8d3e29
0624365c
6fac4f8c
9d2c79c3
125c06c3
235c0484
7f5c0484
37c30021
23974664
402721c3
41c32d35
2a5480c7
0007cf5c
9e0c79c3
42d706c3
25c312c3
01415f5c
466435c3
e3d703b3
365ceaf2
6f8c0624
44cc19c3
0524035c
26641cc3
0624365c
49c36f8c
035c50cc
1cc30644
365c2664
6fac0624
035c50cc
1cc30484
11962664
0f56fc76
00000804
0336f016
61c350c3
0448301c
2010311c
e0cc2c10
0519205c
602644d2
0515305c
00267d0c
0624155c
7cac3664
366405c3
8604201c
2010211c
3364680b
0003351c
401c680e
411c8606
801c2010
811c8606
700b2010
fffd341c
700b700e
60723364
700b700e
fffe341c
700b700e
61723364
0066700e
08959cbc
c007dfe5
201ce794
211c8604
680b2010
fffc341c
28c3680e
341c680b
680efffc
06c37d0c
0624155c
393c3664
64d20014
05c37c4c
60063664
0515355c
0f56c076
00000804
3f36f016
91c3ed96
125c62c3
24370624
893ce8cc
39c3e08c
211c4006
32830800
211c4006
44778000
647762f2
0cb1365c
1c546007
4007402b
32c31954
241c3164
60077fff
323c0a74
04b7ffc0
ae20201c
0011211c
01930d00
ffc0323c
ae20101c
0011111c
24b72c80
40060073
d9c344b7
1000d41c
0044293c
183c4277
2237fff0
01012f5c
50c341f7
023f353c
c01c63b7
193c0000
23770084
0204393c
04576337
02f70172
0024293c
21b342b7
a33c740b
c33c00f4
433c210b
3ac3220b
7b946007
0013a55c
0ac3a085
92dc0007
7d0c000f
241704c3
22973664
6a942007
40074357
3c3c2594
6fd20014
0001831c
375c0494
02330524
0002831c
375c0494
01730564
02537cac
0002c31c
831c1194
05940001
0544375c
01533664
0002831c
375c0494
ff330584
06c37c4c
39c33664
2000341c
600759cc
692c3454
245706c3
59cc3664
080c3a3c
01c321d7
14b40027
22d76037
62062077
60f760b7
00666137
20060177
896c21b7
15c306c3
0300201c
4103211c
60370273
607762d7
00b70206
013700f7
21772066
61b76006
06c3896c
201c15c3
211c1400
60e62010
01534664
06c3692c
36642457
15c30ac3
50bc28c3
3a3c08aa
0f53080c
fff03a3c
78b46027
25d21dc3
03177c0c
36642026
43f7542b
b23ca085
0bc3080c
73540007
20072257
7d0c6394
241704c3
43573664
25944007
00143c3c
831c6fd2
04940001
0524375c
831c0233
04940002
0564375c
7cac0173
c31c0253
11940002
0001831c
375c0594
36640544
831c0153
04940002
0584375c
7c4cff33
366406c3
0dc359cc
1c540007
06c3692c
36642457
3b3c59cc
6037080c
207722d7
60b76046
00f70026
20060137
01b72177
06c3896c
420615c3
4114211c
466460e6
692c0333
1dc306c3
7c0c3664
1dc30dc3
a31c3664
06540002
311c6006
03178000
600602d2
06c36037
404615c3
42bc63d7
3b3c08cd
b580080c
01160153
0b84101c
0000111c
0bc6640c
80563664
32c34397
63b77fe5
00070397
ffef24dc
04d20497
24b72397
393cdb33
60070084
c31c1b94
18940003
0001831c
375c0494
00d30544
0002831c
375c0594
36640584
201c0173
211c0448
680c2010
111c2026
31a30008
1396680f
0f56fc76
00000804
1f36f016
90c3f396
02e4af5c
22771364
836482c3
62373264
60d0a00c
0624655c
2f5cf4cc
42b70121
0544205c
829769ac
425b343c
205c69af
69ac0544
245b383c
305c69af
6dac0544
244b233c
7582301c
2010311c
af5c4c0e
9e100007
425705c3
28c312c3
01014f5c
c66434c3
22f72026
0d91255c
d2dc4007
6257001f
80c743c3
355c0994
6f8c0624
0c8c5ccc
26641ac3
225700b3
420721c3
798921b4
54dc6007
99a9001d
12dc8007
18c3001d
831c24d2
0e940002
0624355c
0f0c6fac
82f78026
0d89155c
d2dc2007
0f4c0008
355c0f73
6fac0624
60260f2c
998907d3
54dc8007
3b69001b
12dc2007
59a9001b
d2dc4007
8257001a
7b8534c3
61873364
355c0db4
28c30624
6fac45f2
60460f4c
6fac0493
80460f6c
225704b3
79e531c3
61e73364
355c0db4
48c30624
6fac85f2
20660f8c
6fac0873
40660fac
825708d3
77e534c3
69e73364
355c0fb4
28c30624
6fac46f2
60860fcc
08b362f7
0fec6fac
82f78086
22570813
321c31c3
3364ff6f
0fb46287
0624355c
86f248c3
035c6fac
20a60404
6fac0373
0424035c
03b340a6
34c38257
ff50321c
63073364
255c18b4
40070d89
38c31454
831c64d2
08940002
0624355c
0f4c6fac
22f720c6
355c0293
6fac0624
40c60f6c
01b342f7
301c0116
311c0b84
6c0c0000
36640a86
60268056
000662f7
1ac37ccc
3a3c3664
60070044
000c14dc
14c38257
37b420c7
0d89255c
400741f7
79e93294
9f2543c3
3f5c81b7
60e700c1
355c0fb4
4f8c0624
9d306fac
125c05c3
235c0484
4f5c0464
34c300e1
39e9c664
5fe521c3
3f5c4177
60a700a1
000999dc
0624255c
435c6bac
6b8c0444
035c5ccc
1ac30644
355c2664
6fac0624
035c5ccc
07730444
31c32257
33647f25
51b460e7
0d89355c
60076137
99e93394
3fe514c3
3f5c20f7
60a70061
355c0fb4
4f8c0624
9d306fac
125c05c3
235c0484
4f5c0444
34c30081
39e9c664
5f2521c3
3f5c40b7
60e70041
255c5d35
6bac0624
0464435c
5ccc6b8c
0644035c
26641ac3
0624355c
5ccc6fac
0464035c
26641ac3
7aa90953
21c32257
359432e4
323c5a49
60070014
62172b94
2d946007
60277a89
063c2a94
101c02c0
111c4b40
fcbc004c
035308b0
22577aa9
32e421c3
5a491c94
0014323c
12946007
60076217
7a891494
11946027
6e6c75cc
02c0063c
4b40101c
004c111c
07f23664
323c10b3
60070024
000812dc
3a2d2006
680c29c3
0007af5c
03c39ef0
13c36257
4f5c28c3
34c30101
8006c664
01411f5c
28c339ed
355c46f2
6f8c0624
02538fec
0001831c
355c0794
6f8c0624
0404435c
831c0133
06940002
0624355c
435c6f8c
7ccc0424
1ac304c3
5a493664
0014323c
75cc6bf2
063c6e6c
101c0340
111c4b40
3664004c
323c00d3
00260044
03c362f2
02b1265c
602645f2
02b5365c
00070073
4bc34654
05c3708c
36642046
19ef30c3
90ec1a0f
040c19c3
5a6913c3
30c34664
63373064
43177b88
34e442c3
1f5c0d54
3b8d0181
03e1255c
7fe532c3
4f5c6077
455c0021
1bc303ed
29c364ac
39ec080c
36644006
70cc4bc3
040c19c3
400639ec
02b33664
42f74026
355cd9b3
6f8c0624
035c5ccc
1ac30644
355c2664
6fac0624
035c5ccc
1ac30484
f0132664
2bc338c4
09c3886c
f88c133c
23c362d7
46646257
01614f5c
7d6c99cd
396905c3
7c6c3664
366405c3
315c19c3
001c06c4
011ceb10
2c4c0009
301c4066
311c0fe4
6cac0000
08745abc
f8760d96
08040f56
ff967016
426441c3
526452c3
04cc204c
200c353c
60264e00
200d233c
62c3678c
c0076383
67cc2494
40072383
343c2094
7580080c
6c006612
343c4c0f
013c0200
7e663a1d
ff7f201c
301ca9d2
311cffff
201cfff3
211cffff
23a3ff7f
343c2083
213c0200
40063b9d
00934037
0096601c
2f5cc037
02c30001
0e560196
00000804
08b8b0bc
00000804
08b8b8bc
00000804
fc961016
31c340c3
60773264
40372364
23c313c3
2d5440a7
13b420a7
40b74006
204713c3
23c36354
04b46047
45944027
605702b3
206713c3
60872d54
02933e94
21c32057
325440e7
20e731c3
23c30a14
14546107
31944127
601702f3
08d3634e
236e2017
3f5c0113
305c0001
07d30225
238e2017
40b74006
3f5c0733
13c30001
08ba0abc
2f5c0633
12c30001
08ba16bc
1f5c0233
20f70001
00612f5c
022d205c
13c332c3
08ba22bc
40170433
4ebc12c3
600608b9
035360b7
31c32057
0010341c
0082101c
600720b7
40571154
51e632c3
60773283
3f5c04c3
13c30021
00013f5c
0cbc23c3
200608b9
2f5c20b7
02c30041
08560496
00000804
fe961016
42c331c3
60373264
23c313c3
18544087
07b42087
602723c3
40670b54
01931c94
13c36017
125420a7
159460c7
234b0073
636b01d3
305c04b3
700e0229
305c0133
700e0221
60776006
238b03d3
4006300e
03334077
31c32017
0010341c
0082101c
60072077
40171054
51e632c3
60373283
00013f5c
f8bc13c3
30c308b8
700e3264
20772006
00212f5c
029602c3
08040856
08b8e2bc
00000804
4e2c604c
21833aa6
4e2f4672
00000804
41c33016
52c34264
204c5264
343c44cc
7580080c
6d006612
341c6c0c
243c8000
6ad20200
2a1d313c
011c0026
30a30001
2b9d313c
313c01b3
40062a1d
0001211c
4026a2f2
343c23a3
213c0200
0c563b9d
00000804
41c31016
22644264
343c004c
303c0200
101c3a1d
111cffff
42f2fffe
13833fc6
0200343c
3b9d103c
08040856
226421c3
323c204c
640500f4
3a1d113c
0080241c
311c6006
42f20001
00066026
62d23183
08040026
326431c3
004c2264
0200133c
303c48d2
40261a1d
0001211c
011332a3
1a1d303c
fffe201c
fffe211c
303c3283
08041b9d
41c33016
52c34264
204c5264
343c44cc
7580080c
6d006612
341c6c0c
243c8000
6ad20200
2a1d313c
011c0806
30a30040
2b9d313c
313c01b3
40062a1d
0040211c
4806a2f2
343c23a3
213c0200
0c563b9d
00000804
51c33016
804c5364
0404345c
345c7672
531c0407
09940400
201c2006
211cc9d0
66a60011
08bc6cbc
5aa6722c
353c3283
722f41ac
08040c56
684c404c
31833706
680c684f
680f6092
680f6046
00000804
204c7016
6092640c
4046640f
640c440f
0002341c
a1467df2
610fa74f
676f612f
23c3806c
601c7100
611c8000
cc0f0040
ac4fa026
231c4805
f5940300
301c84cf
311c0100
6c2c2021
0010341c
662c63d2
40ec662f
8006a14c
a8ef0373
680f6026
601c682c
368380ff
610c682f
410f63f2
612c0093
4c0f6cec
68ec412f
cc0fc006
36c3c3ab
63ae6025
a1854405
305c8025
6ecb0b24
e21443e4
211c4806
215c0040
315c0407
501c0404
511cfffe
3583fffe
0407315c
0147601c
4026c44f
0e56440f
00000804
301c3016
311c0100
6c0c2021
00ff341c
0100201c
2021211c
644f6d00
0e64415c
315c84af
0cac0b24
4ecb04cf
acac4512
654f6a80
04ef846f
00ff201c
01c3474e
08b976bc
0c560006
00000804
604c21c3
025432e4
08040013
32c343cb
63ce6025
00000804
326431c3
233c204c
313c0110
78722a1d
2b9d313c
00000804
326431c3
233c204c
313c0110
77722a1d
2b9d313c
00000804
313c404c
7872c80c
602668af
0804634e
ff96f016
c409a04c
f4cc8429
200c343c
60264f00
200d033c
20c3778c
40072383
57cc4394
328330c3
3e946007
080c363c
66126e00
44498f80
0c944027
6709050b
211c4006
63d24000
f00c233c
812c303c
050b01f3
44ac4ad2
311c6006
42f22000
303c32c3
009381ac
800c303c
700f6f72
343c8409
653c0200
64293a1d
211c4006
63f200c0
00c0201c
02462449
004662f2
313c26a3
23a3000d
0200343c
3b9d253c
40374006
201c0093
40370095
00013f5c
019603c3
08040f56
72c3f016
626461c3
50cc804c
380c363c
533c6d00
700c0280
700f6d72
15c307c3
b0bc4106
700c08cb
2000341c
700c75d2
700f6d92
36236026
0f56736f
00000804
fc963016
a04c40c3
63d2600c
200f2006
341c762c
60070100
762c1c94
2004133c
25d220f7
245c4046
00b30215
00613f5c
0215345c
20372006
0211245c
60064077
00463f5c
22a604c3
32c34006
08bbeabc
233c762c
40070804
734b1194
0080331c
73eb0d94
4037734e
2f5c4077
04c30046
32c32266
08bbeabc
20460073
0496334e
08040c56
434bfd96
201c43ee
434e0080
60376006
3f5c6077
22860046
eabc23c3
039608bb
00000804
fb963016
804c50c3
20372006
40062077
00462f5c
40062206
eabc32c3
70ac08bb
ffff101c
01ff111c
70af3183
736f736c
73ef73ec
3ff2338c
53af5fe6
02d32137
3f5c05c3
13c30081
e2bc4006
05c308b8
00812f5c
402612c3
08b8e2bc
13c36117
20f72025
00612f5c
355c4137
21170219
32e421c3
722ce6b4
0100341c
11546007
740f6026
374e2066
40374006
60064077
00463f5c
220605c3
eabc32c3
009308bb
76bc05c3
059608b9
08040c56
2026fc96
105c2037
20770e64
1f5c2026
12c30046
600623c3
08d1babc
326430c3
64d260f7
0094301c
1f5c60f7
01c30061
08040496
404c1016
88cc228c
31542007
6baf6046
341c6bac
7df20002
604600f3
6bac6baf
0002341c
6bcc7df2
0002341c
440c77f2
23837c06
640f6026
63f2610c
0093210f
6cec612c
212f2c0f
200664ec
23ab2c0f
602531c3
12c363ae
ea944007
0800343c
205c428f
20260407
4c6f2c4f
08040856
30c3ff96
40a63264
64d24037
00ff201c
3f5c4037
03c30001
08040196
326430c3
7f5233c4
400603c3
2021211c
080402a3
326430c3
7f5233c4
201c03c3
211c0100
02a32021
00000804
08ba22bc
00000804
f6961016
01814f5c
4f5c8077
1f5c01a1
3f5c0045
2f5c004d
2f5c00c6
2f5c0021
81f70055
104b243c
3f5c4037
3f5c0001
1f3c0105
2abc0080
0a9608ba
08040856
fc967016
c21760f7
13648257
01433f5c
220760b7
22071754
27d203b4
228706f3
22a71a54
04d33394
1f5c8037
1f5c0041
12c30025
00613f5c
36c323c3
08c2a2bc
305c04b3
80370b44
00411f5c
00251f5c
01338e2c
0b44305c
1f5c8037
1f5c0041
8e0c0025
3f5c12c3
23c30061
466436c3
803701b3
00411f5c
00251f5c
3f5c12c3
23c30061
ccbc36c3
000608bc
0e560496
00000804
fd963016
026451c3
22640077
301c4037
8c0c0b00
0e64045c
0300101c
08cb9cbc
0b24345c
4ecb0cac
02c7123c
08cb9cbc
345c60a6
1f5c020d
145c0001
2f5c021d
02c30021
d8bc14c3
30c308b9
201c3264
40b7008d
940f63f2
3f5c60b7
03c30041
0c560396
00000804
08b96abc
00000804
2006fc96
0001111c
105c2037
28050e64
20262077
00461f5c
23c312c3
babc6026
30c308d1
60f73264
301c64d2
60f70093
00611f5c
049601c3
00000804
060c301c
4130311c
40066c0c
0010211c
6dd23283
feb0303c
09b46027
313c0006
331c808c
04544105
00530026
08040006
10c3f016
c197e157
536452c3
2f5c3264
405c00e1
60070b44
49d21794
0b24305c
65f26ccc
15c371ec
02533664
0b89315c
039460a7
0053912c
01c3910c
26c315c3
466437c3
602700b3
714c0394
0f563664
00000804
00213f5c
0215305c
00000804
4e2c604c
4e2f4672
00000804
08e4305c
4d0d5f46
00000804
205c1016
313c0b24
880c280c
40806e00
325c2dcb
13e405e1
64060634
4110311c
8c0f8206
08040856
0136f016
70c3fc96
0b24005c
280c323c
cd00400c
504b41c3
a0061010
600770cb
375c1294
001c0211
60470200
08060254
341d2006
62f23200
013c2026
00f70016
00615f5c
38ac788c
18cc2037
5f5c0077
07c30046
babc18c3
70cb08d1
60078105
aef2db94
38ac788c
58cc2037
00264077
00460f5c
18c307c3
babc25c3
049608d1
0f568076
00000804
fd963016
428c50c3
880c0273
60376046
0e64355c
0080321c
40b76077
202605c3
60464006
08d468bc
7c0624c3
40072383
0396ed94
08040c56
fe967016
660660c3
4105311c
0c0e0226
265cc077
365c0b64
60a70b89
301c0e94
311cc200
690f0001
525ca006
525c0125
0106012d
0135025c
0140301c
2021311c
233c6c0c
40370014
4007a057
355c6054
0cac0b24
153caecb
9cbc02c7
605708cb
0480033c
9cbc2c06
605708cb
0d0f0006
0d2f6057
20066057
40572fae
0b24325c
a8cfacac
215c2057
6acb0b24
08ac6512
654f6c00
2cac6057
60572c6f
4cef4ccc
8d4c6057
00062cec
84ef0333
640f6026
690c4057
290f63f2
692c0093
2c0f6cec
2d2f6057
a00664ec
4057ac0f
35c3abab
6bae6025
81852405
40570025
0b24325c
03e46ecb
0046e314
05ed025c
345c8057
ae4c0b44
200606c3
345c40e6
56640b81
335c6057
20260b24
0d732c8f
0b44355c
06c38e4c
40c62086
0b81355c
2f5c4664
02c30001
00401f3c
34bc40c6
30c308bc
62d23264
40570013
0b89325c
0f946087
ca1c001c
0011011c
08c7025c
101c6057
111cca80
135c0011
01d308e7
ca08301c
0011311c
08c7325c
501c6057
511cca3c
535c0011
605708e7
0f80033c
08c4135c
b0bc4246
405708cb
0f80323c
08c7325c
235c6057
435c08e4
033c08e4
12c31200
b0bc502b
405708cb
1200323c
08e7325c
001c6057
011cca30
035c0011
60570867
cabc101c
0011111c
0887135c
323c4057
325c0d80
005708a7
402620c6
08b7e6bc
0e560296
00000804
305cff96
133c08e4
21c3039e
00bf241c
1f5c4037
2c0d0001
400620c6
08b7e6bc
08040196
fd96f016
51c340c3
40b72264
0653205c
705c5012
cb800663
0649205c
365442c7
795442e7
c4dc42a7
02c30008
8abc16c3
000708bc
0008e4dc
b2dca007
345c0008
70120653
0663145c
145c4c80
20870673
208710b4
e80c0594
0547745c
20470113
480b0394
48090053
0547245c
0a80243c
200604c3
0673345c
08bc6cbc
200604c3
32c34006
08bb50bc
02c30c93
8abc16c3
000708bc
a0075e94
345c2154
70120653
0663545c
245c4e80
045c0567
345c05a7
60870673
243c06b4
20260b00
05a7145c
200604c3
0673345c
08bb50bc
200604c3
32c34006
08bc6cbc
345c0793
600705a4
545c3854
345c05a7
60870673
345c0794
545c0564
ac0f0584
245c0593
445c0564
80770584
03946047
0473880e
00211f5c
03f3280d
1d542007
40062006
50bc32c3
04c308bb
40062006
6cbc32c3
345c08bc
6dec0b44
145c04c3
36640653
205c0153
82170b44
88cc8037
00415f5c
466425c3
0f560396
00000804
ff961016
200740c3
68091c54
06546027
21c32006
08b7e2bc
682b0293
08896037
213c3000
341c681e
23e400ff
3f5c0454
640d0001
200604c3
32c34006
08bc6cbc
08560196
00000804
21c32006
08b7e2bc
00000804
f9967016
305c60c3
61b708e4
42dc2007
682b0010
141c13c3
131cff00
72dc0300
131c0009
09d40300
0100131c
131c0f54
64dc0200
0253000e
0600131c
000ab2dc
0700131c
000dd4dc
465c1593
686b08c4
09dc6227
6246000d
365c19b3
20b70211
03546047
60b76806
0b89365c
4d946087
0f5c6197
00370041
00011f5c
61972ecd
a832a097
0f5ca077
0eed0021
1f5c6197
2fad0001
5f5c6197
afcd0021
0f5c6197
035c0001
61970125
00211f5c
012d135c
5f5c6197
535c0001
6197015d
00210f5c
0165035c
1f5c6197
135c0001
61970195
00215f5c
019d535c
0f5c6197
035c0001
619701cd
00211f5c
01d5135c
486ba197
6c2b6197
34e442c3
619703b4
06c38c2b
25c32006
01d334c3
0e9460a7
686b8197
482b4197
03b423e4
6c2b6197
200606c3
6cbc24c3
365c08bc
8e4c0b44
200606c3
365c40e6
46640b81
0b44365c
06c38e4c
40c620a6
0b81365c
0c134664
0ff4133c
02f420e7
365c2106
133c0e04
64091a1d
886b03c3
236423c3
336434c3
023523e4
50c304c3
a9675364
00130235
1720463c
25c304c3
08cbb0bc
200606c3
35c324c3
465c0693
686b0864
2c356127
05536146
0211365c
0200001c
604700f7
68060354
365c60f7
5f5c0884
a1370061
00810f5c
365c0ecd
20d70884
21772832
00a15f5c
365caeed
0f5c0884
0fad0081
0884365c
00a11f5c
465c2fcd
686b0884
02356767
06c36786
24c32006
08bc6cbc
06c300f3
21c32006
08b7e2bc
06c300f3
40062006
50bc32c3
079608bb
08040e56
50c37016
200742c3
c8092454
0794c047
08e4305c
6c894889
067423e4
21c32006
08b7e2bc
20a602d3
08a4205c
08b862bc
08a4255c
6027706b
36c30235
200605c3
08bc6cbc
200605c3
32c34006
08bb50bc
08040e56
ff967016
61c340c3
202652c3
00202f3c
08b862bc
00131f5c
04c327d2
21c32006
08b7e2bc
c00702d3
54891454
321c32c3
518000d0
346b31c3
602622d2
200604c3
08bc6cbc
200604c3
32c34006
08bb50bc
0e560196
00000804
fe963016
52c340c3
44542007
20372849
04f42027
21c32006
2f3c0473
60170060
21946007
62bc2026
3f5c08b8
60270033
04c312b4
60172086
e6bc23c3
04c308b7
40262026
08b7e6bc
2f5c04c3
12c30001
03b34017
3f5c04c3
13c30001
e2bc23c3
031308b7
62bc2086
3f5c08b8
54490033
055432e4
208604c3
08b7e6bc
202604c3
e6bc4006
04c308b7
40062006
6cbc32c3
029608bc
08040c56
ff961016
200740c3
20861854
00202f3c
08b862bc
08a4345c
00112f5c
04c34c0d
245c2006
602608a4
08bc6cbc
200604c3
32c34006
08bb50bc
08560196
00000804
fc963016
52c340c3
65542007
40774809
404744d2
07b35694
6027742b
60470454
01d33394
2f3c20c6
62bc00e0
2f5c08b8
41720073
00762f5c
20c604c3
748907f3
65f26037
0211305c
03546047
073304c3
2f3c2026
62bc00e0
3f5c08b8
60470073
60260bb4
06a6345c
32c3544b
ff00341c
06b6345c
04c30533
00013f5c
23c313c3
08b7e2bc
2f5c0633
12c30021
ff1332c3
4007542b
54891694
341c32c3
6472008f
3f5c60b7
13c30041
00e02f3c
08b862bc
2f5c04c3
12c30041
e6bc4026
009308b7
21c32006
04c3fbd3
40062006
6cbc32c3
015308bc
06a3305c
305c67d2
20e606b3
e6bc23c3
049608b7
08040c56
fd96f016
61c340c3
7f3c52c3
202600a0
62bc27c3
3f5c08b8
60270053
c0073fb4
74094254
64d26037
38946047
742b0333
10946027
20c604c3
62bc27c3
3f5c08b8
23c30053
fffd241c
00562f5c
20c604c3
04c30393
00012f5c
21c312c3
d42b0453
1c94c007
32c35489
008f341c
60776472
3f5c04c3
13c30021
62bc27c3
04c308b8
00212f5c
26c312c3
08b7e6bc
200604c3
32c34006
08bc6cbc
04c300d3
21c32006
08b7e2bc
0f560396
00000804
fb963016
503c40c3
20070c30
68094954
0081331c
331c0c54
15540082
0080331c
20c63b94
62bc25c3
053308b8
41806889
01403f3c
0681225c
fc7e233c
23c32006
04336086
31c3284b
008f341c
60376472
00012f5c
2f3c12c3
62bc0120
3f5c08b8
60770091
00211f5c
061d145c
00932f5c
40b74832
00413f5c
0625345c
200604c3
604625c3
08bc6cbc
200604c3
32c34006
08bb50bc
200600b3
e2bc21c3
059608b7
08040c56
fe967016
305c50c3
601c0211
60470200
c8060254
436446c3
3f5c6046
40260005
00252f5c
12c305c3
600624c3
08bbcabc
3f5c6046
40260005
00252f5c
12c305c3
31c324c3
08bbcabc
3f5c6046
40260005
00252f5c
13c305c3
600624c3
08bbcabc
3f5c6046
40260005
00252f5c
13c305c3
602624c3
08bbcabc
3f5c6046
40260005
00252f5c
206605c3
600624c3
08bbcabc
3f5c6046
40260005
00252f5c
206605c3
602624c3
08bbcabc
0b44355c
05c36dac
366416c3
0b44355c
05c38e4c
40e62006
0b81355c
355c4664
40260b24
02964c8f
08040e56
40c31016
48492cd2
e6bc2066
04c308b7
40062006
6cbc32c3
00b308bc
40262026
08b7e6bc
0b24345c
64f26c8c
1cbc04c3
085608c2
00000804
0336f016
50c3fd96
93c361c3
40b72264
0c80703c
0b64405c
200625d2
86bc27c3
855c08ba
831c0b89
5d940005
0641355c
241c23c3
4077001f
55944027
0649355c
06546427
25546447
48946407
c0070233
05c34a54
243c2006
60e60200
08bc6cbc
200605c3
32c34006
08bb50bc
c0070793
05c33a54
243c2006
355c0200
50bc0673
05c308bb
40062006
6cbc32c3
057308bc
2954c007
0651255c
3f5c05c3
13c30021
08b7e6bc
200605c3
32c34006
08bc6cbc
0653255c
341c32c3
60070002
355c1454
40570b24
355c4c8f
8e4c0b44
18c305c3
355c40c6
46640b81
05c300d3
21c32006
08b7e2bc
0641255c
341c32c3
64070060
68076954
60077254
355c7d94
60e70649
60e73d54
60670fb4
60672754
600706b4
60271754
03536f94
245460a7
6a9460c7
614704f3
61473d54
610706b4
61272d54
06136194
3a546167
5c946187
05c307b3
27c316c3
08c1cabc
05c30b53
27c316c3
08c174bc
05c30a93
27c316c3
08c0febc
05c309d3
27c316c3
08c286bc
05c30913
27c316c3
08bf2ebc
05c30853
27c316c3
08bf28bc
05c30793
27c316c3
08c0debc
05c306d3
27c316c3
08c092bc
05c30613
27c316c3
08c066bc
05c30553
27c316c3
08bf04bc
05c30493
27c316c3
08c03cbc
355c03d3
8cec0b44
16c305c3
00413f5c
37c323c3
02734664
0b44355c
40374297
05c38cac
3f5c16c3
23c30041
466439c3
05c300d3
21c32006
08b7e2bc
c0760396
08040f56
00000804
005c7016
205c05c4
313c0724
880c280c
95ebae00
0187343c
0704405c
68abce00
1b9431e4
04946027
0ba4405c
405c0073
542b0bc4
7fe532c3
742e3364
71806412
0c2c584c
26642006
6412742b
40067180
742b4c2f
ee946007
08040e56
0014313c
201c69d2
211c00ac
680c4140
60073164
4606fdd4
4105211c
3364680b
680e6172
662c204c
66727792
2606662f
4105111c
341c680b
7ad20040
341c640b
640effd9
0b24305c
4e4e4006
00000804
605c7016
265c05c4
20470704
313c20b4
a9800187
06c3748c
554b2006
30c33664
43c33264
1e546007
06c3742c
36642006
000740c3
01161794
0b84301c
0000311c
001c6c0c
366400d4
01938056
301c0116
311c0b84
6c0c0000
00d5001c
80563664
04c38006
08040e56
05c4305c
494c4d6c
266403c3
00000804
0f36f016
b0c3f996
805ca3c3
605c05c4
401c0b64
f1200200
315c18c3
6c4c0764
74dc6007
515c0008
55090ea4
75292264
233c3264
7549412c
233c3264
7569812c
c12c333c
15806185
27c31ac3
08cbb0bc
22645509
32647529
412c233c
32647549
812c233c
333c7569
7d80c12c
0ff4133c
55092137
00812f5c
233c550d
40f7420b
1f5c5529
352d0061
440b133c
554920b7
00412f5c
233c554d
4077c08c
3f5c7569
756d0021
22645509
32647529
412c233c
32647549
812c233c
333c7569
6067c12c
453c3435
550900c0
75292264
233c3264
7549412c
333c3264
5569812c
14c30ac3
c1ac223c
08cbb0bc
22645509
32647529
412c233c
32647549
812c233c
733c7569
04c3c12c
cc20101c
0011111c
44bc4086
01640892
235c38c3
303c0764
33c40b0d
60257f32
00b3684f
1ac30bc3
143324c3
315c18c3
4c4c0764
19944027
37c35811
784e3364
78eb586e
236423c3
34dc4007
780c0009
784b784f
78ee3364
586e584e
0166644c
a2bc2c0c
10b30872
915c18c3
29c30ba4
6007682c
3ac33994
656cac0c
053c6cec
36641b0b
326430c3
602661b7
31232197
437223c3
0ba0301c
0000311c
21832c0b
41b742f2
323c4197
18c30187
0704115c
001c8c80
011c0bb4
15c30000
088bbabc
00c12f5c
39c35b8d
78af6c2c
fff4253c
66ec18c3
68802f0c
500b78cf
68a0302b
4006792e
3b895a0d
0187313c
225c28c3
8d000704
18ac592b
0bb472e4
27c31ac3
08cbb0bc
6f8078ac
392b78af
047367a0
b0bc1ac3
5a0908cb
602532c3
1f5c6037
21770001
00a12f5c
31c35a0d
19c36412
6c2c6580
592b78af
3ac303c3
5d202d00
08cbb0bc
7d20592b
6c8038ac
300b78af
6fa06880
78cc792e
78cf6fa0
706c64f2
366408c3
1ac30bc3
0200201c
08c69ebc
f0760796
08040f56
02c330c3
135c26f2
a2bc0b81
02930872
12542027
10542047
0e542067
06942087
0b81135c
0872e8bc
20a700f3
135c0594
16bc0b81
08040873
0b00301c
00e66c0c
0b81135c
087300bc
00000804
40c37016
05c4505c
0b24605c
0361155c
62942007
211c4606
680b4105
351c3364
680e0024
6a2c404c
31833aa6
6a2f7772
6c2c744c
0b946087
301c0116
311c0b84
6c0c0000
00d1001c
80563664
0111365c
01166bf2
0b84301c
0000311c
001c6c0c
366400d2
20068056
0115165c
10c30006
087348bc
11540007
6c2c744c
0d946047
0edc301c
0000311c
67f26c0c
0f14301c
0000311c
6cd26c0c
1388001c
08959cbc
0b44345c
04c36c8c
36642006
345c02b3
535c0b24
a0470131
00260b94
0b81145c
0872d0bc
145c05c3
d0bc0b81
345c0872
20260b24
0e562e4e
00000804
305c3016
6ceb0b64
305c69d2
8e4c0b44
41662006
0b81305c
0c564664
00000804
fc961016
01004f3c
ffde143c
0b24305c
233c6c0c
688c0200
203728ac
207728cc
2f5c4026
14c30046
babc4026
049608d1
08040856
fd967016
405c51c3
304c0b64
11542007
0b24305c
233c6c0c
682c0200
c037c84c
c077c86c
2f5c4026
25c30046
08d1babc
70ee6006
706b70ce
60273364
700c0994
704b704f
70ee3364
504e4006
0396506e
08040e56
ff963016
105c51c3
64eb0b64
8e247fd2
64cbf524
444c3364
60376d22
602564cb
64ce3364
7fe564eb
64ee3364
64f264eb
34bc15c3
343c08c6
62d24004
3f5cf324
03c30001
0c560196
00000804
fd967016
536452c3
636463c3
1054a007
0b24305c
233c6c0c
688c0200
803788ac
807788cc
00466f5c
babc25c3
039608d1
08040e56
fd963016
0b24305c
433c6c0c
702c0200
a037b04c
a077b06c
4f5c8026
babc0046
039608d1
08040c56
1264fd96
60062264
60776037
68bc60b7
039608d4
00000804
08b79ebc
00000804
0080301c
4040311c
0100201c
301c4c0e
311c0db0
40060000
620c4d0d
20866c2c
08043664
0080301c
4040311c
0800201c
301c4c0e
311c0db0
40060000
101c4d6d
111c0b54
f0bc0000
08040873
0080301c
4040311c
0400201c
301c4c0e
311c0db0
40060000
301c4d4d
311c0fe4
2cac0000
0873f0bc
00000804
0fe4301c
0000311c
f0bc2ccc
08040873
0fe4301c
0000311c
f0bc2c8c
08040873
0fe4301c
0000311c
f0bc2cec
08040873
0f36f016
70c3fe96
0080201c
4040211c
313c080b
2486080c
4080111c
6c0b6c80
13e33364
20771083
00215f5c
c006a80e
4040611c
0db0b01c
0000b11c
0daca01c
0000a11c
0b84901c
0000911c
0001801c
05c304b3
08ce0cbc
436440c3
0067343c
782cd980
0204233c
45f24037
00011f5c
2e213bc3
680c2ac3
4a1d333c
07c364d2
00f33664
19c30116
0f66640c
80563664
400d383c
358333e3
a00753c3
0296db94
0f56f076
00000804
16bc2066
080408c7
16bc2046
080408c7
16bc2026
080408c7
16bc2006
080408c7
0736f016
650670c3
4110311c
313c4c0c
2486080c
4080111c
6c0b6c80
33e33364
41dc323c
536453c3
a01cc026
a11c0024
901c4110
911c0dac
801c0000
811c0b84
03f30000
0cbc05c3
40c308ce
343c4364
363cff80
2ac3300d
19c3680f
333c640c
64d24a1d
366407c3
011600f3
680c28c3
36640f46
363c8056
33e3400d
53c33583
e194a007
0f56e076
00000804
7abc2066
080408c7
7abc2046
080408c7
7abc2026
080408c7
7abc2006
080408c7
0336f016
61c340c3
23942007
311c6406
6c0b4080
001c3364
011cdd00
80270000
001c0e54
011cee00
89d20000
bb00001c
0000011c
03548047
7700001c
400613c3
0810211c
63127100
32646c0b
041303a3
01c32006
1c94c027
311c6446
6c0b4080
47863364
4080211c
123c480b
343c81ac
0086180c
4080011c
4c0b6c00
01662364
1020011c
62127000
033c6c0b
50e3812c
901c5183
911c0f38
801c0000
811c0b84
e0260000
05c303d3
08ce0cbc
303c40c3
c0270100
30c30254
303c09c3
67d23a1d
0bb4001c
0000011c
00f33664
28c30116
0f26680c
80563664
400d373c
538333e3
e294a007
0f56c076
00000804
20260066
08c7d0bc
00000804
20260046
08c7d0bc
00000804
10c30026
08c7d0bc
00000804
20260006
08c7d0bc
00000804
20060066
08c7d0bc
00000804
20060046
08c7d0bc
00000804
20060026
08c7d0bc
00000804
10c30006
08c7d0bc
00000804
08fd3abc
00000804
60c3f016
42c351c3
f524ee24
78bc0f86
053c08cc
143c0340
40260a1d
600d323c
343c31a3
25230b9d
311c6406
4c0f4110
82bc0f86
373c08cc
62d24004
0f56f324
00000804
60c3f016
52c341c3
f524ee24
78bc0f86
243c08cc
153c0340
60262a1d
33e33623
353c3183
0f862b9d
08cc82bc
4004373c
f32462d2
08040f56
60c3f016
52c341c3
f524ee24
78bc0f86
243c08cc
153c0300
60262a1d
33e33623
353c3183
0f862b9d
08cc82bc
4004373c
f32462d2
08040f56
60c3f016
42c351c3
f524ee24
78bc0f86
053c08cc
143c0300
40260a1d
600d323c
343c31a3
25230b9d
311c6406
4c0f4110
82bc0f86
373c08cc
62d24004
0f56f324
00000804
0136f016
41c380c3
53c372c3
011c0006
64001044
4c0c6212
31236026
111c2486
640f4110
5fe75fe5
0f86fd94
08cc78bc
0300243c
2a1d153c
0340343c
3a1d453c
153c4183
34e32a1d
353c3183
0f862b9d
08cc82bc
1a548007
501cc026
511c0b84
04c30000
08ce0cbc
000d263c
428322e3
0a1d373c
08c364d2
00d33664
740c0116
36640ec6
80078056
8076ed94
08040f56
0fe4301c
0000311c
20666d0c
0900233c
08c8f6bc
00000804
0fe4301c
0000311c
20466d0c
0600233c
08c8f6bc
00000804
0fe4301c
0000311c
20266d0c
0300233c
08c8f6bc
00000804
0fe4301c
0000311c
20066d0c
f6bc23c3
080408c8
804c1016
0306600c
1341135c
0872b8bc
345c6026
345c0195
7ef201a1
08040856
4046600c
1345235c
20460306
0872a2bc
00000804
8e241016
31e3f524
3283402c
64f2602f
70bc00ab
343c0895
62d24004
0856f324
00000804
40c33016
f524ae24
66d2602c
70bc00ab
60060895
353c702f
62d24004
0c56f324
00000804
f5240c16
00040004
20c30004
301c2364
311c0244
4c0e2020
311c6086
40864105
301c4c0e
311c0844
41e62200
30564c0f
08040013
a06c3016
311c6186
6c0c4140
0ae1205c
011c0006
42f24000
4fe602c3
ffff211c
313c3283
30a351ac
211c4186
680f4140
fff0213c
6506948c
210d033c
466415c3
08040c56
40c33016
700c52c3
0001341c
702c6bd2
5e7223c3
311c6186
4c0f4140
05c3648c
aee73664
63860735
4105311c
53724c0c
638600d3
4105311c
53924c0c
300c4c0f
0084313c
504c67d2
4008301c
4128311c
313c4c0f
67d20104
301c506c
311c400c
4c0f4128
301c508c
311c4000
4c0f4128
08040c56
0bb4301c
0000311c
48cc4e0c
266403c3
00000804
0bb4301c
0000311c
2c4c4e2c
03c3482c
26642b05
00000804
0bb4301c
0000311c
2c4c4e2c
03c3482c
0098121c
08042664
ff96f016
605c50c3
e20c06e4
612c804c
36646dcc
6dac752c
366405c3
341c706c
60070001
01061954
08881ebc
0fe4301c
0000311c
00066d4c
9000011c
36643fe6
6c6c752c
36640fc3
582c6017
782f6d20
6d00580c
7c2c784f
202605c3
355c3664
6fd20c44
0128301c
4130311c
03ff201c
301c4c0f
311c0088
201c4080
4c0f1fff
0f560196
00000804
1f36f016
90c3fc96
600c6070
c48c8e50
333c782c
3364650b
1bc36037
202687cc
600641c6
70c34664
4eac39c3
17c4335c
3f866065
125c3183
4c8004a4
0200301c
a0c32d20
801ca284
20070001
1bc32b94
29c364cc
2026080c
a0c33664
0010183c
073c20f7
383c1f9d
6312fff0
782c5d80
650b333c
063e123c
680e65a0
180c383c
782c5d80
650b333c
275c68ce
32c30293
375c6025
3f5c0296
83c30061
101c8264
782c0200
51c37432
023553e4
984c53c3
0007af5c
333c782c
3264120b
a0b76077
011c0006
1cc31000
101c201c
0000211c
8cbc34c3
784c08a4
784f6e80
a00c253c
6d20782c
2006782f
400643c3
fff0211c
80074283
1bc3ab94
0404315c
17c309c3
04c33664
f8760496
08040f56
0336f016
60c3ff96
82c371c3
021793c3
2587b80c
06d20794
05c30037
088ababc
746c0453
8fcc0037
17c305c3
39c328c3
40c34664
17c4355c
5f866065
41803283
333c680c
680f232b
19c0063c
420612c3
08cbb0bc
345c6006
79cc0286
06c36cac
366414c3
c0760196
08040f56
40c31016
f5240e24
0edc201c
0000211c
6025680c
684c680f
282f63f2
2c2f0053
0edc301c
0000311c
60062c4f
303c642f
62d24004
704cf324
2c0c00c6
0872a2bc
08040856
21c31016
27e730c3
80061535
8c2f8c0f
8c6f8c4f
8caf8c8f
8cef8ccf
8d2f8d0f
8d6f8d4f
8daf8d8f
8def8dcf
38056805
123cfd73
780603f4
01002383
31c320c3
093561e7
880f8006
884f882f
4205886f
fef37e05
00f4213c
0304313c
40670180
80060635
027f403c
ff535f85
08040856
50c37016
0034613c
5f8641c3
14c34283
08cb64bc
1600c8d2
40066006
602541a1
fc9463e4
08040e56
0f36f016
a1c390c3
32c362c3
31833f86
838480c3
f1804ac3
bc0003c4
840018c3
74300193
346c544c
084f353c
7031700f
306f504f
82050205
f4741e27
38c34006
3c008c00
a5010093
4085b161
7fa76800
263cfb74
48d20034
19c37920
4ac30580
5ebc3180
f0760891
08040f56
08cbb0bc
00000804
50c37016
02c341c3
35a26006
12e451a2
00460334
12e40133
00260335
602500b3
f49403e4
0e560006
00000804
0084301c
4140311c
600f6c0c
00000804
0114301c
4130311c
133c6c0c
301c104b
311c8218
001c2404
011c3333
0c0f0033
8208201c
2404211c
0006680c
0180011c
680f30a3
14942007
680c4085
111c2006
31a300a0
4085680f
0006680c
0002011c
7bd23083
8200301c
2404311c
20270313
201c1894
211c820c
680c2404
011c0006
30a30140
4085680f
2006680c
0001111c
7bd23183
8214301c
2404311c
04130c0c
13942047
820c201c
2404211c
0006680c
0340011c
680f30a3
680c4085
111c2006
31830001
fcf37bd2
301c0116
311c0b84
6c0c0000
00b5001c
80563664
203c0006
301c488c
311c0080
4c0f4140
00000804
8000201c
1040211c
233c6100
680c100c
08047ff2
8000201c
1040211c
62126100
4c0f4006
00000804
3f36f016
00f7fc96
42c381c3
4007d3c3
301c7054
311c456c
6c0c4114
080cc23c
a026e006
0056323c
0b0d333c
933c7fe5
0ad3f88c
40d71984
0d91625c
233c38c3
323c161d
c3f24d8b
450b323c
621219a4
4000201c
4114211c
0c0c6d00
139480a7
c7006bc3
c045c077
4006c0b7
233c63d7
6057671d
402523c3
808c303c
363cc3d7
0473271d
c8d24680
633c63d7
a6c3259d
ffc0a41c
63d700f3
259d633c
a41ca6c3
c3d7fff0
271da63c
40774680
808c603c
62c3a6c3
323c43d7
23c3659d
af5ca2a3
63d70047
671da33c
6700c017
023c43d7
20a5371d
af1414e4
e0258c84
7de4b600
b73c0834
353c0057
6037fff0
fe732006
fc760496
08040f56
0511105c
301c29d2
311c0448
4c0c2010
4c0f4072
201c0173
211c0448
680c2010
111c2026
31a30008
0804680f
0511105c
301c29d2
311c0448
4c0c2010
4c0f4092
201c0193
211c0448
680c2010
fffe101c
fff7111c
680f3183
00000804
800c1016
6dac60cc
70cc3664
04c36cac
08563664
00000804
1f36f016
51c3c0c3
83c392c3
b23ce297
8006080c
fff0633c
a364a7c3
253c0853
3cc3161d
0d91335c
323c6ed2
62124d8b
4000001c
4114011c
001c6c00
011cffff
01b3003f
450b323c
001c6212
011c4000
6c004114
ffff001c
000f011c
4c0f2083
19e42045
46e4dd14
5b840554
6007742b
eed21794
135446e4
0ac38025
0415e007
0df2142b
0bd2140b
08959cbc
34c30113
333c3603
33c40b0d
91807f32
8025a085
033448e4
fbd32006
0f56f876
00000804
800c1016
6c4c60cc
345c3664
6dac0544
fe00201c
0001211c
01463283
03c662d2
08959cbc
6d8c70cc
366404c3
08040856
40c37016
52c361c3
6ad241a6
60274286
43860754
04546047
04946067
42e442c6
01160b14
0b84301c
0000311c
001c6c0c
36640091
343c8056
1580100c
6cd2600c
301c0116
311c0b84
6c0c0000
0092001c
80563664
c00f0053
08040e56
40c33016
61a651c3
62864ad2
07544027
40476386
40670454
62c60494
0a1443e4
301c0116
311c0b84
6c0c0000
366401a6
343c8056
9580100c
6bf2700c
301c0116
311c0b84
6c0c0000
0090001c
80563664
500f4006
08040c56
333c30c3
333c080d
03c30b8d
00000804
0336f016
70c3ff96
00f0a04c
0001901c
76ac07d3
0cbc03c3
40c308ce
78bc0ee6
56ac08cc
400d693c
328336e3
0ee676af
08cc82bc
0280343c
3a1d453c
70695029
0001341c
1d946007
32647069
60376072
00011f5c
7069306d
0010341c
323c69f2
5580300c
384e123c
31a336c3
55ec680f
393c3009
32a3100d
74ac75ef
74af6025
69ec28c3
366407c3
708d6006
600776ac
0473c194
03c3762c
08ce0cbc
0ee640c3
08cc78bc
363c362c
23e3400d
318332c3
766c762f
138312c3
768c366f
568f2383
82bc0ee6
343c08cc
18c30280
07c344ec
3a1d153c
00532664
762cc026
db946007
c0760196
08040f56
70c3f016
4006804c
524e520e
704f6006
53c364c3
0504165c
25d2a025
6c8c7e0c
366407c3
a087c085
704cf694
05946047
6c0c7d2c
366407c3
375c6006
0f5604c5
00000804
804c1016
0361305c
62cc6bd2
36646c8c
0026303c
0b0d333c
7f3233c4
60260053
085671cf
00000804
404c3016
0644405c
00270449
a54b0894
aa0b35c3
6a0e35a3
0193084f
0a940047
6027684c
084f0254
30c3058b
30a30a4b
684c6a4e
03946027
00539009
88ef9029
08040c56
0336f016
50c3fd96
04a4105c
68942007
311c6646
00264105
60450c0e
355c4c0b
4c0e0684
311c6786
4c0b4105
0684355c
76ec4c2e
455c0e70
04c30664
683c21c3
763c108c
0653100c
301c92c3
311c01fa
93842020
6c0939c3
92c36037
01fc301c
2020311c
39c39384
60776c09
301c92c3
311c01fe
93842020
6c0939c3
92c360b7
01f8301c
2020311c
39c39384
70a16c09
00013f5c
ffed305c
00213f5c
fff5305c
00413f5c
fffd305c
41052085
17e40085
363ccc94
001c180c
011c0200
4c002020
48c33080
0100001c
1010011c
61127000
423c00b3
413c011f
23e400df
4026fb94
04a7255c
c0760396
08040f56
ff963016
5f5c81cc
a0370083
1264908c
32642264
01964664
08040c56
40c37016
62c34364
343c6364
201c100c
211c0f38
ad000000
6cd2740c
301c0116
311c0b84
6c0c0000
008c001c
80563664
340f0053
0d3583e7
100c363c
211c45c6
2d004080
fe00243c
32236026
02b3640f
0104343c
180c263c
60c668d2
4080311c
441c4980
00b3ffef
311c6046
49804080
34236026
680e3364
0e5605c3
00000804
03641016
303c2364
401c100c
411c0f38
2e000000
0104303c
323c6ad2
8086180c
4080411c
041c4e00
00f3ffef
411c8006
6a000810
180c233c
30236026
680e3364
64d2640c
640f6006
01160173
0b84301c
0000311c
001c6c0c
3664008c
00068056
08040856
50c37016
62c35364
353c6364
201c100c
211c0dac
080c0000
700c8c00
01166cd2
0b84301c
0000311c
001c6c0c
36640094
00538056
363c300f
4486080c
4080211c
640b2d00
40263364
22e32523
640e3283
0e5604c3
00000804
600f6006
080c313c
111c2486
0c804080
6026200b
200d233c
32c321a3
600e3364
08040006
0136f016
70c381c3
62c37364
301c6364
311c0fe4
ad0c0000
60c645c3
1254c007
0300453c
c0276106
453c0d54
60860600
0854c047
0900453c
c0676146
60060354
336443c3
0b1473e4
301c0116
311c0b84
6c0c0000
009a001c
80563664
100c373c
680c5180
01166cd2
0b84301c
0000311c
001c6c0c
36640093
00538056
0f860811
08cc78bc
0340163c
1a1d353c
27234026
353c32a3
0f861b9d
08cc82bc
0f568076
00000804
40c33016
0084201c
4140211c
082c280c
31e4680c
300ffc14
0c56102f
00000804
0336f016
82c371c3
440c43c3
202848d2
43e46500
68a004d4
181543e4
313c10c3
d1a0018f
61126048
ffe0533c
60684006
04f463e4
25e40045
9c0f0714
2c296500
340d58c3
40450073
c076fe73
08040f56
1f36f016
a2c371c3
2f5c83c3
244b0141
341c31c3
6007000f
80863a94
53c303c3
c2c35c6b
0002c21c
0001901c
b43c05b3
3ac30010
68494c00
c8297012
41ac363c
c4221ac3
31a316c3
363cc869
3563c1ac
c40918c3
293c16c3
5fe5100d
2bc33283
271d373c
821c68c3
363c0001
5580009f
190c323c
03c36180
523c0364
343c0074
43c30020
c4e44364
0b13d315
4d946027
61127c6b
936493c3
305c46f2
6fac0624
01f3cecc
231cc006
0b5400ff
301c0116
311c0b84
6c0c0000
36640c06
c0068056
0006a086
921c40c3
b01c0002
05530001
44221ac3
2e2238c3
0f352107
800c323c
41ac323c
223c32a3
3b3cc1ac
7fe5100d
303c2383
00f30020
100d3b3c
23837fe5
0010303c
036403c3
080c353c
3a227d80
2c0c2123
4c0f21a3
0020353c
536453c3
95e48025
0153d615
301c0116
311c0b84
6c0c0000
36640be6
f8768056
08040f56
0736f016
80c3f996
51c3a2c3
93c35064
4f5c9364
600c01e0
0624735c
3370083c
0b33c006
fff8105c
0241275c
341c32c3
62d20002
28c38068
335c680c
602703d1
c0672a94
313c0bb4
5f890030
6e806d20
61b76e00
00c13f5c
c1670773
5f8909b4
6e806520
61776e00
00a13f5c
5f890633
6ad239c3
ffd0313c
6e806d20
61376e00
00812f5c
652003b3
6e006e80
3f5c60f7
03d30061
09b4c0e7
65205f89
6e006e80
3f5c60b7
02930041
39c35f89
313c6bd2
6d20ffd0
6e006e80
2f5c6077
400d0021
65200113
6e006e80
3f5c6037
600d0001
0205c025
a7146ae4
325c28c3
4ca904c4
28c347d2
335c686c
08c30704
07963664
0f56e076
00000804
0f36f016
af5c81c3
e2970124
936493c3
01636f5c
505c804c
210c0b24
64ec28d2
610f6c0c
45946007
0873612f
323c0013
351c800c
00938080
800c323c
642f6772
0c5164ec
644c0451
1000321c
293c646f
303c0120
a0062a1d
103c64f2
a0262b9d
01e0393c
3a1d203c
3b9d103c
280f42d2
1794a007
0ac3738c
00070383
700c2994
700f6e72
2ac373cc
700c2383
4000341c
700c77d2
700f6e92
1a944007
00733c4f
40063c4f
07c35c6f
08b9febc
02135391
b3c363ab
ffffb21c
01d6b05c
b3c376eb
0001b21c
0176b55c
b794c027
0006f633
0f56f076
00000804
3f36f016
b0c3d396
0b24a05c
21b7204c
2027276c
61060a94
a0066037
00255f5c
600625c3
08c2a2bc
03ec0197
21970237
400607ef
239743b7
62171364
32dc6007
20a7001f
60260eb4
833c0397
4217000d
91c38283
62b76006
a00758c3
3b331394
30c30397
40266145
300d823c
83836217
a00758c3
001ce2dc
ffa0313c
936493c3
38e342b7
21c32217
42372383
080c393c
2e80a297
00c0213c
303c0ac3
60252a1d
2b9d303c
d364d1c3
01203d3c
153c5bc3
01973a1d
3d3c40cc
c3c3300c
8006c284
02978377
261c20c3
41770001
fff0393c
f88c033c
013702a3
05c4a297
32d300f7
00070117
642c1754
0080341c
10546007
6027640c
0018e2dc
6c2c640c
0080341c
74dc6007
642c0018
642f6792
62972ff3
642c6bd2
0080341c
642c67f2
8000341c
a02663d2
642ca377
7c0b233c
640c4337
3583bc06
642c61f7
0684233c
427702c3
341c4ad2
67d20040
4c6c3cc3
328330e3
606f0cc3
6c4c64ec
40d762f7
600732c4
931c3754
34940001
100c343c
0010743c
00070357
2f3c2754
69800b40
ff47135c
09c06f3c
0373a006
059454e4
0ac32026
0316105c
00078f5c
0027cf5c
40b7580c
20260bc3
3dc321c3
08d468bc
3ac30006
0316035c
163c2006
a025027f
e51457e4
5f3c2613
75800b40
ff47135c
60071c13
931c3754
34940002
100c343c
0010743c
40074357
5f3c2754
75800b40
fe87135c
08406f3c
0373a006
059454e4
1ac34026
0326215c
00078f5c
0027cf5c
60b7780c
20460bc3
3dc34026
08d468bc
0ac32006
0326105c
263c4006
a025027f
e51457e4
5f3c1f13
75800b40
fe87135c
60071513
931c3754
34940003
100c343c
0010743c
40074357
5f3c2754
75800b40
fdc7135c
06c06f3c
0373a006
059454e4
1ac34026
0336215c
00078f5c
0027cf5c
60b7780c
20660bc3
3dc34026
08d468bc
0ac32006
0336105c
263c4006
a025027f
e51457e4
5f3c1813
75800b40
fdc7135c
60070e13
931c3754
34940004
100c343c
0010743c
40074357
5f3c2754
75800b40
fd07135c
05406f3c
0373a006
059454e4
1ac34026
0346215c
00078f5c
0027cf5c
60b7780c
20860bc3
3dc34026
08d468bc
0ac32006
0346105c
263c4006
a025027f
e51457e4
5f3c1113
75800b40
fd07135c
60070713
931c3854
35940005
100c343c
0010743c
40074357
5f3c2754
75800b40
fc47135c
03c06f3c
0373a006
059454e4
1ac34026
0356215c
00078f5c
0027cf5c
60b7780c
20a60bc3
3dc34026
08d468bc
0ac32006
0356105c
263c4006
a025027f
e51457e4
5f3c0a13
75800b40
fc47135c
027347c3
00070117
8f5c1054
cf5c0007
20b70027
19c30bc3
23c36297
68bc3dc3
59c308d4
1d54a007
04f202d7
22d22157
43570013
21d745f2
60076157
a2d72154
0317a037
1f5c0077
1f5c0121
0bc30045
29c32006
01415f5c
a2bc35c3
01f308bc
00370317
01211f5c
00251f5c
19c30bc3
01413f5c
62d723c3
08c2a2bc
200721d7
ffe6a4dc
05c3a397
03b70025
e4dc0187
0073ffe0
f9338006
fc762d96
08040f56
301c7016
ac0c0b00
982cd44c
3483784c
21546007
343c982f
64d20014
26bc05c3
343c08d2
64d20404
fabc05c3
343c08ba
64d20044
a6bc05c3
343c08ba
64d20024
04bc05c3
343c08ba
60071004
05c3df54
08bae8bc
08040e56
0736f016
c21750c3
01249f5c
13648297
a364a2c3
836483c3
005ce04c
42eb0b24
7fe532c3
c00762ee
3a3c1694
4c80200c
633c6026
313c200d
4ac3080c
83c37180
5ccc8364
300c383c
928493c3
0120383c
3a1d453c
04942027
0313205c
204702b3
205c0494
02130323
04942067
0333205c
20870173
205c0494
00d30343
20a74006
205c0394
80070353
300c5754
10831c06
341c702c
60070080
dfaf1054
06c37fac
1df20383
dfaf00d3
06c37fac
1df20383
06c37fcc
18f20383
700f6026
63f2750c
0093950f
6cec752c
952f8c0f
800670ec
17ab8c0f
602530c3
2ef277ae
0120383c
3b9d153c
01e0383c
3b9d153c
29c36026
286f684f
44f20433
80074ac3
383c1d94
153c0120
642c3b9d
0080341c
14546007
7fccdf8f
038306c3
7f8c0ff2
238326c3
7fcc5df2
438346c3
09c387f2
806f204f
08b9febc
0006df8f
0f56e076
00000804
3f36f016
50c3ff96
c3c362c3
05c4705c
0b24a05c
280c313c
000c0ac3
5c0c8c00
81c34037
0ac38364
0056805c
4cd228c3
0a5481e4
301c0116
311c0b84
6c0c0000
36640226
11cb8056
7fe530c3
945c71ce
19c300f3
d75c24f2
00730ba4
0bc4d75c
0187393c
275cb3c3
b2840704
155c00e6
00bc0b81
3bc30873
62e44c0b
1ac31794
6025642c
500b642f
01164bd2
0b84301c
0000311c
001c6c0c
36640086
0bc38056
0cc3604c
36642006
cb200c33
331c700b
0e3501ff
01ff631c
01160bb4
0b84301c
0000311c
001c6c0c
36640086
5cc38056
6007700b
0ac31b94
0056805c
815c1bc3
5cc30013
340b5884
fff4313c
42ac0017
04c4025c
700e6c00
45f229c3
6dac7d6c
366407c3
600668a4
845c702e
383c0013
0dc3200c
ac2f6180
302bcc4f
602531c3
700b702e
0b3436e4
301c0116
311c0b84
6c0c0000
0086001c
80563664
6320100b
236423c3
4007500e
383c1194
60a70010
641206b4
61800dc3
4c2f4c4f
646c1bc3
366407c3
2ac36006
019668ae
0f56fc76
00000804
3f36f016
d0c3fc96
0b00201c
2e24a80c
f52420f7
0b24355c
75c38c0c
8405c026
00f3845c
0187383c
115c1dc3
4c800704
6007696b
90302854
50707050
0003925c
355c03b3
6d8c0b44
18c305c3
10c33664
19540007
0b00201c
bf5c680c
af5c0007
40260027
00462f5c
29c303c3
babc3cc3
31cb08d1
602531c3
51cb71ce
05e9375c
e01423e4
e025c025
6b8c2dc3
61e413c3
00e6c735
0b81155c
0872d0bc
32c340d7
0400341c
f32462d2
fc760496
08040f56
1f36f016
62ec80c3
405c8e70
74c30664
56c3c006
108cac3c
100cba3c
175c03f3
075cffe9
975cfff1
301cfff9
311c01f8
55802020
680e7322
01fa201c
2020211c
2c0e7500
75004045
001c0c0e
011c01fe
74002020
0006935c
e085c085
6be4a105
3300df94
180c3a3c
0200401c
2020411c
0cc34e00
0100401c
1010411c
61126200
013c00b3
023c009f
23e4015f
08c3fb94
0684105c
6686440b
4105311c
442b4c0e
4c0e6105
311c6646
40464105
600c4c0e
0d23235c
0246301c
2020311c
f8764c0e
08040f56
0f36f016
80c3ff96
4006a04c
00062f5c
00162f5c
6429f60c
0a946027
012c301c
4130311c
60376c0c
447223c3
40060153
07946067
012c301c
4130311c
40374c0c
315c18c3
69d20c44
008c301c
4080311c
641ccc0c
06f31407
00a8301c
4140311c
633c6c0c
05f300c4
0cbc07c3
40c308ce
0280303c
3a1d253c
31c3294b
0203341c
c00763d2
298b1094
0014313c
39c363d2
313c6af2
63d22004
25f219c3
341c6869
6cf20002
6a2c28c3
08c36c4c
366414c3
3bc304c3
b4bc2c6c
3a3c0873
33e3400d
01937383
0fe4b01c
0000b11c
0b0d323c
933c33c4
a01cf88c
e0070001
18c3c694
0c44315c
68f247c3
00a8301c
4140311c
433c6c0c
770c0204
12546007
033c76cc
340c0010
0872a2bc
6b2c28c3
08946087
76cc87d2
0010033c
d0bc340c
01960872
0f56f076
00000804
00000001
00080010
003c0103
00070107
0004011e
00050121
00000001
00080010
003c0103
00090107
0005011e
00030121
00000001
00080010
00500103
00060107
0003011e
00040121
00000001
00080010
00200103
00030107
0002011e
00050121
00000001
00080010
00300103
00060107
0004011e
00070121
00000001
00760110
04000002
040200ff
00070005
6630000f
0f090018
9231001a
4ddf001b
4537001d
0f120024
00a00029
3000002a
00010036
0347003a
8411003b
5f63004b
00370059
ffff00be
000000bf
07770306
03330307
7bde030a
0200030b
71ff030c
00700311
e0c10314
29200352
0000011b
01360162
00e60163
08440800
00c80808
00c80809
d5df080a
c00e080b
000c011d
117d0150
080a0119
00000129
000b016f
00100160
00450f00
104b0133
014c014e
003c0123
0caa0106
50180149
a0940026
e8000325
0b200165
0200012f
01220162
00d80163
01000079
fcb800c4
1c040116
40000021
0000007c
000a0300
80000f01
00000001
00340110
b7f40364
9d260365
ee100366
37be0367
3cfc0368
05570369
c0cc036a
9723036b
e83c036c
386b036d
906d037c
c74a037d
2414037e
3175037f
3e530380
05ca0381
96210382
bd300383
200d0384
35c30385
c000036e
40000386
4000037a
0a09006f
0001006e
00300012
00000001
00300110
00c80808
00a00029
0f120024
000a0322
903d0134
00800011
3d510017
9ee60045
05940055
c5c1005d
fcb800c4
666a0009
3d510017
0064001e
0064001f
9233003f
c6100040
006f0041
00530042
9ee60045
08660049
05940055
00000015
80000020
00000001
00040111
4ef57000
4c3f0808
403fbc00
0000000a
00000001
00020111
403fbc00
00000190
00000001
001f0111
5581fe00
55c09020
4cc00000
40a04000
40400000
42000000
4d300000
4c3f0820
4d74c410
4de00000
4e2a1000
4f400000
4ef57000
4f150008
483e8000
48800006
54400000
54800000
54c00000
00000100
54c0f7b0
54204c00
00000064
485e6120
41724c00
568207b0
447a0000
44280000
44d0c120
4510c120
45c12000
00000001
00020111
40000000
55800000
00000001
00030031
403fbc00
5581fe00
000000c8
00000001
00050111
40a04000
54c17bd0
485e2120
0000000a
445a0000
00000001
00010111
44780000
00000001
00150111
40a04000
445a0000
41c00000
4c3f0820
48800006
54c17bd0
485e2120
0000000a
5628b100
5628b180
0000003c
48840206
00000014
48860306
0000001e
48870386
00000032
4c3f0808
48870382
41e93900
0000000a
00000001
00020111
403f7c00
00000190
00000002
00020110
01000f01
001d0111
5588be00
55c08020
4cc00000
40a04000
40400000
42000000
4d300000
4c3f0820
4d7501a0
4dda0000
4e2a1000
4f6d0020
4edbb00c
4f150000
483e8000
48800006
54400000
54800000
54c0f7b0
54204c00
00000064
485e6120
568207b0
44bd0000
442b8400
4570c600
45b0c600
45c12000
41724800
00000001
00020111
40000000
55800000
00000001
00030031
403f7c00
5588be00
000000c8
00000001
00820110
fffc0302
40040303
60000003
8214000d
00800011
002e00aa
003c0102
003c0104
003c0105
002a0108
0030010a
002c010b
002c010c
0014010e
298a0111
38880112
50c80113
380a0114
01e40115
1c1c011c
0016011f
1a240120
00070121
00140122
00320125
00240126
00200127
00600128
903d0134
9030013b
0e0d0146
01ea014b
0801014c
000a015d
1510015e
5021015f
00d20312
00610301
0524030f
72c00323
37a90324
3da0034f
01000319
0000031a
0000031b
0000031c
0100031d
0000031e
100a0322
00000348
39eb0f03
04670f05
00a30f07
00f20f09
0ef00f0b
00130f0d
ff580f04
0f800f06
00580f08
0f6c0f0a
00de0f0c
0ff90f0e
25c20f0f
00d80f10
00000f02
00000001
00340111
4d7501a0
4dda0000
503b9800
50433000
50800000
50c0b700
483e0000
44780000
503b8000
4ef57000
568207a0
40d60000
41998000
5114a420
68020000
68421000
68822000
68c40000
69041000
69442000
69860000
69c61000
6a062000
6a463000
6a864000
6ac82000
6b083000
6b484000
6b885000
6bc86000
6c087000
6c488000
6c889000
6cc8a000
6d08b000
6d48c000
6d88d000
6dc8e000
6e08f000
6e490000
6e891000
6ec92000
6f093000
6f494000
6f895000
6fc96000
41c00000
4c3f0808
48870382
0000000a
41e93900
40a14000
00000002
00f40110
01000f01
fffc0302
40040303
60010003
8214000d
00c00011
00e00035
86800046
00010058
002e00aa
003c0102
003c0104
003c0105
00280108
002c010a
002c010b
002c010c
000c010e
298a0111
3a880112
52c80113
380a0114
01e40115
1b1b011c
0016011f
1a260120
00160122
00500125
00200126
00200127
01e00128
000a012a
000a012b
0100012f
903d0134
9030013b
1e0d0146
01ea014b
0001014c
0006015d
01c2015b
1510015e
3021015f
00d20312
00610301
72c00323
37a90324
3da0034f
01000319
0000031a
0000031b
0000031c
0100031d
0000031e
100a0322
00000348
36440f03
07ff0f05
00a10f07
0d5e0f09
0f0b0f0b
00900f0d
f9df0f04
04c70f06
00960f08
0a320f0a
07c10f0c
0ede0f0e
25c20f0f
00d80f10
00000f02
02603008
07e03009
0404300a
0040300b
0000300c
0002300d
0000300e
0000300f
02763010
03763011
00063012
00403013
00003014
00023015
00003016
00003017
02763018
06ae3019
0000301a
0040301b
0000301c
00a2301d
0000301e
0000301f
02603048
00003049
0000304a
0040304b
0000304c
0002304d
0000304e
0000304f
02763050
00003051
00003052
00403053
00003054
00023055
00003056
00003057
02763058
00003059
0000305a
0040305b
0000305c
00a2305d
0000305e
0000305f
14370022
040a0023
0f120024
002c0111
523b9800
52424c80
52a00000
52c0b700
483e0000
44bc0000
523b8000
4edbb00c
568207a0
40f20000
41a1c000
53294948
68020000
68421000
68822000
68c23000
69024000
69442000
69843000
69c44000
6a062000
6a463000
6a864000
6ac82000
6b083000
6b484000
6b885000
6bc86000
6c087000
6c488000
6c889000
6cc8a000
6d08b000
6d48c000
6d88d000
6dc8e000
6e08f000
6e490000
6e891000
6ec92000
6f093000
6f494000
6f895000
6fc96000
00000002
00020030
386100ab
00030031
485e6120
48786120
40a54000
00000002
00100030
486100ab
4531001d
000b010e
0005015d
1510015e
000d0160
1a240120
0030010a
00030031
485ea120
4878a120
40a54000
00000002
00020030
386100ab
00030031
485e2120
48782120
40a54000
00000002
00020030
386100ab
00040031
54c17bdc
485e2120
48782120
40a54000
00000001
00040111
d6400000
ca800000
ca000000
ca400000
00000001
00030111
ce800000
d5000000
cd400000
00000001
00050011
5589fe00
00000064
56c00000
56e00000
0000012c
00000001
00000111
403fbc00
00000001
00030111
4f6d0020
4f150000
4570c600
00000001
00030111
4f6d0000
4f00000c
4570c698
00000001
00010111
449d0000
00000001
00010111
44bc0000
00000001
00130111
40a04000
41c00000
4c3f0820
48800006
54c17bd0
485e2120
5628b100
5628b180
0000003c
48840206
00000014
48860306
0000001e
48870386
00000032
4c3f0808
48870382
0000000a
41e93900
00000001
00000111
403f7c00
00000001
00050111
4e2a1000
4f150008
54c0f7b0
44d0c120
49820000
00000001
00050111
4e001000
4f150004
54c0d7b0
44d10120
49a00000
00000001
00050111
4e001000
4f100000
54c0d7b0
44d101b0
49a00000
00000001
00050111
4e2a1000
4edbb00c
54c0f7b0
45c12000
49820000
00000001
00050111
4e2a1000
4edbb00c
54c0d7b0
45c12000
49820000
00000001
00080111
4e001000
4f100000
4f6d0000
4edbb000
54c0d7b0
45710010
45c12010
49820000
00000001
00020111
5114a420
40d60000
00000001
00020111
51086210
40d60000
00000001
00020111
51002000
00000000
000040d2
00000001
00020111
5310c850
40f20000
00000001
00020111
c6100002
00005310
000040f2
00000001
00020111
53104000
40f20000
1919191a
00000019
00010020
000d0009
0061001a
00a10081
00e100c1
00620062
00a20082
00e200c2
00c300a3
008500e3
00c500a5
00e600e5
00e800e7
00ea00e9
00ef00ec
00f400f4
00f400f4
00f400f4
000000f4
0004001d
000d000b
000b0019
0019000d
000d000b
000b0019
0019000d
00060006
00060006
00260007
00460045
00660047
00860067
00880087
00a80089
00e800a9
00ea00e9
00ed00eb
00f000ee
00f200f2
00f200f2
000600f2
00060006
00070006
00450026
00470046
00670066
00870086
00890088
00a900a8
00e900e8
00eb00ea
00ee00ed
00f200f0
00f200f2
00f200f2
00060006
00060006
00260007
00460045
00660047
00860067
00880087
00a80089
00e800a9
00ea00e9
00ed00eb
00f000ee
00f200f2
00f200f2
000600f2
00060006
00070006
00450026
00470046
00670066
00870086
00890088
00a900a8
00e900e8
00eb00ea
00ee00ed
00f200f0
00f200f2
00f200f2
0e0e0e0e
0a0a0a0a
0a0a0a0a
0a0a0a0a
0a0a0a0a
0e0e0e0e
0a0a0a0a
0a0a0a0a
0a0a0a0a
0a0a0a0a
0e0e0e0e
0a0a0a0a
0a0a0a0a
0a0a0a0a
0a0a0a0a
0e0e0e0e
0a0a0a0a
0a0a0a0a
0a0a0a0a
0a0a0a0a
0c0c0c0b
0a0a0a0a
0a0a0a0a
0a0a0a0a
090a0a0a
02020202
02020200
020202ff
02020202
fdff0002
03030300
03030300
03030303
00000003
03030300
03030300
03030303
00000003
03030300
03030300
03030303
00000003
03030300
03030300
03030303
00000003
03030300
03030300
03030303
00000003
03030300
03030300
03030303
00000003
03030300
03030300
03030303
00000003
03030300
03030300
03030303
00000003
03030300
03030300
03030303
00000003
09090906
09090905
09090909
04050609
09090906
09090905
09090909
04050609
09090905
09090904
09090909
03040509
09090905
09090904
09090909
03040509
fdfdfdfb
fdfdfdfa
fdfdfdfd
f9fafbfd
fdfdfdfb
fdfdfdfa
fdfdfdfd
f9fafbfd
fcfcfcfa
fcfcfcf9
fcfcfcfc
f8f9fafc
fdfdfdfa
fdfdfdf9
fdfdfdfd
f8f9fafd
00000001
00010111
48800002
00000001
00010111
4d74c410
00000001
00010111
4d7501a0
00000001
00c00110
00000170
00040171
00080172
000c0173
00100174
00140175
00180176
001c0177
00200178
00240179
0028017a
002c017b
0030017c
0034017d
0038017e
003c017f
00400180
00440181
00480182
004c0183
00500184
00540185
00580186
005c0187
00600188
00640189
0068018a
006c018b
0070018c
0074018d
0078018e
007c018f
00020190
00060191
000a0192
000e0193
00120194
00160195
001a0196
001e0197
00220198
00260199
002a019a
002e019b
0032019c
0036019d
003a019e
003e019f
004201a0
004601a1
004a01a2
004e01a3
005201a4
005601a5
005a01a6
005e01a7
006201a8
006601a9
006a01aa
006e01ab
007201ac
007601ad
007a01ae
007e01af
000301b0
000701b1
000b01b2
000f01b3
001301b4
001701b5
001b01b6
001f01b7
002301b8
002701b9
002b01ba
002f01bb
003301bc
003701bd
003b01be
003f01bf
004301c0
004701c1
004b01c2
004f01c3
005301c4
005701c5
005701c6
005701c7
005701c8
005701c9
005701ca
005701cb
005701cc
005701cd
005701ce
005701cf
00000001
00c00110
04100170
04110171
04120172
04200173
04210174
04220175
04300176
04310177
04320178
04400179
0441017a
0442017b
0443017c
0444017d
0445017e
0446017f
04470180
04480181
04490182
044a0183
044b0184
044b0185
044b0186
044b0187
044b0188
044b0189
044b018a
044b018b
044b018c
044b018d
044b018e
044b018f
02100190
02110191
02120192
02200193
02210194
02220195
02300196
02310197
02320198
02400199
0241019a
0242019b
0243019c
0244019d
0245019e
0246019f
024701a0
024801a1
024901a2
024a01a3
024b01a4
024b01a5
024b01a6
024b01a7
024b01a8
024b01a9
024b01aa
024b01ab
024b01ac
024b01ad
024b01ae
024b01af
001001b0
001101b1
001201b2
002001b3
002101b4
002201b5
003001b6
003101b7
003201b8
004001b9
004101ba
004201bb
004301bc
004401bd
004501be
004601bf
004701c0
004801c1
004901c2
004a01c3
004b01c4
004b01c5
004b01c6
004b01c7
004b01c8
004b01c9
004b01ca
004b01cb
004b01cc
004b01cd
004b01ce
004b01cf
00000001
00400110
00000002
fffc0302
40040303
32c00323
20100c03
0c8a0106
002a0108
21860111
06080112
00d00113
08080114
94c90115
0014011f
00100122
00100125
00240126
00180127
00600128
0001014c
5f0e015e
5009015f
04000c05
000c011d
000b016f
01000319
0000031a
0000031b
0000031c
0100031d
0000031e
000a0322
00600301
00000001
000d0111
4d74c410
4de00000
503b9800
50438400
50800000
50c0b700
40a14000
483e0000
44780000
503b8000
4ef57000
568207a0
5114a420
00000001
00a60110
8214000d
00d20312
00540102
00500104
00500105
0050010a
0050010b
0050010c
0010010e
060a0112
9cc90115
00140119
1d1d011c
12280120
00020131
903c0134
00b0013b
0001014c
0006015d
ca4b0c04
0b800c06
16700c07
15020c08
1d4c001c
00000c40
eaaa0c41
00010c42
eb000c43
04000c05
00050c49
00000c4b
0200030d
3e20034f
0bff0507
0bff0506
0bff0509
0bff0508
0c1a050b
0c4e050a
0c3e050d
0c83050c
0c4c050f
0b2e050e
0b050511
0ac00510
0ab30513
0ab20512
0ab8051c
0aa5051b
0a28051e
0a06051d
0a540520
0aa5051f
0af30522
0bb80521
0c4e0524
0d200523
0e140526
00000525
00000528
00000527
00000514
00000515
00000516
00000517
00000518
00000519
0000051a
00000529
0000052a
0000052b
0000052c
0000052d
0000052e
0000052f
00000c53
00000c54
00000c55
00000c56
00000c4f
1fa40c4e
1f480c4d
1eec0c4c
00000001
00320111
41998000
5114a420
40a14000
485e2120
4c3f0820
48800006
54400000
54800000
54c1fffc
540afc00
00000064
48782120
68020000
68421000
68822000
68c40000
69041000
69442000
69860000
69c61000
6a062000
6a463000
6a864000
6ac82000
6b083000
6b484000
6b885000
6bc86000
6c087000
6c488000
6c889000
6cc8a000
6d08b000
6d48c000
6d88d000
6dc8e000
6e08f000
6e490000
6e891000
6ec92000
6f093000
6f494000
6f895000
6fc96000
41c00000
4c3f0808
48870382
0000000a
41e93900
4d74c410
00000001
00010111
54301c00
00000001
00010111
54351c00
00000001
00010111
54207c00
00000001
00010111
54207c00
00000002
000a0110
0fde0c58
00320c57
02100c50
60100c5e
09000c51
00010111
54207c00
00000002
000a0110
97020c08
60080c48
00800c4a
00000c5e
01000146
00010111
54191c00
00000001
00010111
543f1c00
00000002
000a0110
97010c08
af260c48
01000c4a
00030c5e
00000146
00010111
5419fc00
00000001
00640110
8214000d
0fd20312
00200102
001c0104
001c0105
008a0106
0018010a
0014010b
0014010c
0010010e
04880112
30500113
1d1d011c
0c0c0120
01ff012a
01020131
903c0134
0070013b
01e2014b
0001014c
0006015d
0a450c04
0b800c06
02700c07
000c011d
000b016f
90000c08
00000c40
df9f0c41
00010c42
0e000c43
04000c05
79df0c48
00000c49
00800c4a
00000c4b
8a0f0c52
00000c50
00000c51
00000c5e
0200030d
28000323
3e20034f
00000c65
00000503
0b00003e
5009015f
21800111
08040140
01000146
00000001
00310111
41998000
40a14000
485e2120
4c3f0820
48800006
54400000
54800000
54c1fffc
54351c00
00000064
48782120
68020000
68421000
68822000
68c40000
69041000
69442000
69860000
69c61000
6a062000
6a463000
6a864000
6ac82000
6b083000
6b484000
6b885000
6bc86000
6c087000
6c488000
6c889000
6cc8a000
6d08b000
6d48c000
6d88d000
6dc8e000
6e08f000
6e490000
6e891000
6ec92000
6f093000
6f494000
6f895000
6fc96000
41c00000
4c3f0808
48870382
0000000a
41e93900
4d74c410
00000002
00020110
90e00c08
00010111
5419fc00
00000002
00040110
0c8a0106
90020c08
00010111
5419fc00
00000001
00060110
0030013b
d9990c41
00040c65
00000001
00060110
0030013b
d6960c41
00080c65
00000001
001c0110
00400125
060f0112
02b0013b
00100c09
903d0134
e4640c41
69df0c48
00080c49
00900c4a
5a00001c
c1000146
9a0f0c52
66000c65
00000503
00000001
00140110
00100125
04880112
0070013b
903c0134
de9e0c41
1d4c001c
8a0f0c52
00000c65
00000c6a
00000503
00000001
002e0110
0214000d
0fd20312
00300102
00300104
00300105
0030010a
0030010b
0030010c
0014010e
1616011c
161a0120
00100c09
903d0134
01b0013b
000d015d
c2f00c04
a6800c06
07100c07
00f10c08
00400c20
36540c21
00000c22
3e20034f
00000001
00300111
419dc000
40a14000
485e2120
4c3f0820
48800006
54400000
54800000
54c17bdc
5411fc00
00000064
48782120
68020000
68421000
68822000
68c40000
69041000
69442000
69860000
69c61000
6a062000
6a463000
6a864000
6ac82000
6b083000
6b484000
6b885000
6bc86000
6c087000
6c488000
6c889000
6cc8a000
6d08b000
6d48c000
6d88d000
6dc8e000
6e08f000
6e490000
6e891000
6ec92000
6f093000
6f494000
6f895000
6fc96000
41c00000
4c3f0808
48870382
0000000a
41e93900
00000001
00040031
54c1fffc
485e2120
48782120
40a54000
00000001
00040031
54c17bdc
485e2120
48782120
40a54000
00000001
00010031
40a54000
00000001
00010111
4d74c410
522b5441
00000000
4a3205fd
512f7874
1481eb10
b8c953ca
0a601907
00000002
7d8f90ad
81fe115f
20e9ce42
213b333b
0923bb58
332c7f8c
647ede6c
00000066
00000c8c
00001920
000025b0
00003240
00004b64
00006488
00007118
00007dac
00001918
00003234
00004b50
0000646c
000096a8
0000c8e0
0000e1fc
0000fb18
0000259c
00004b3c
000070e0
00009680
0000e1c0
0000fffc
0000fffc
0000fffc
0000321c
00006438
00009658
0000c878
0000fffc
0000fffc
0000fffc
0000fffc
00000df4
00001be8
000029e0
000037d8
000053c4
00006fb4
00007dac
00008ba0
00001be4
000037cc
000053b4
00006f98
0000a768
0000df38
0000fb20
0000fffc
000029cc
000053a0
00007d70
0000a740
0000fae4
0000fffc
0000fffc
0000fffc
000037b0
00006f64
0000a71c
0000ded0
0000fffc
0000fffc
0000fffc
0000fffc
00001a18
00003430
00004e4c
00006864
00009c9c
0000d0d0
0000eaec
0000fffc
00003424
0000684c
00009c74
0000d098
0000fffc
0000fffc
0000fffc
0000fffc
00004e24
00009c48
0000ea70
0000fffc
0000fffc
0000fffc
0000fffc
0000fffc
00006814
0000d02c
0000fffc
0000fffc
0000fffc
0000fffc
0000fffc
0000fffc
00001cfc
000039fc
00005700
00007400
0000ae00
0000e804
0000fffc
0000fffc
000039f0
000073e4
0000add8
0000e7cc
0000fffc
0000fffc
0000fffc
0000fffc
000056d8
0000adb0
0000fffc
0000fffc
0000fffc
0000fffc
0000fffc
0000fffc
000073b0
0000e760
0000fffc
0000fffc
0000fffc
0000fffc
0000fffc
0000fffc
0036001a
006c0034
00a2004e
00d80068
0144009c
01b000d0
01e600ea
021c0104
00020001
000b000b
060c1830
09122436
0036001a
00ea0075
006c0034
01d400ea
00a2004e
02be015f
00d80068
03a801d4
0144009c
057c02be
01b000d0
075003a8
01e600ea
083a041d
021c0104
09240492
02880138
0af8057c
02d00000
0c300618
00000000
00000000
aaaaaa00
aaaaaaaa
eeeeeeaa
eeeeeeee
fffffeee
ffffffff
ffffffff
dfbf7fff
fdfbf7ef
dfbf7efc
fdfbf7ef
0000007e
02000112
40000002
91161618
02010002
00000100
02000112
40ffffff
91161618
02010002
00000106
0200060a
40ffffff
00000001
00430209
c0000102
00040932
02020100
24050001
05011000
00010124
02022404
00062405
82050701
0b004003
00010409
00000a02
81050700
00020002
02010507
00000200
003c0209
c0040101
00040996
ffff0600
050700ff
00400281
01050700
00004002
02820507
07000200
00020205
05070002
02000283
03050700
00020002
003c0709
c0040101
00040996
ffff0200
050700ff
02000281
01050700
00004002
02820507
07000040
40020205
05070000
00400283
03050700
00004002
00000007
04090304
0052032c
00640065
00690070
0065006e
00530020
00670069
0061006e
0073006c
0020002c
006e0049
002e0063
00570338
00720069
006c0065
00730065
00200073
00530055
00200042
0065004e
00770074
0072006f
0020006b
006f004d
00750064
0065006c
00570340
00720069
006c0065
00730065
00200073
00530055
002d0042
00440043
00200043
0065004e
00770074
0072006f
0020006b
006f004d
00750064
0065006c
0042030a
00540045
00000041
00230308
00320030
005f0308
00310041
0030031a
00300030
00300030
00300030
00300030
00300030
00000031
0059031e
0075006f
00200072
0061006e
0065006d
00680020
00720065
00000065
00420322
00440041
00530020
00520054
004e0049
00200047
006e0049
00650064
00000078
522b5441
00000000
42c33016
702c442c
0a9423e4
240c402f
12e4500c
200f0334
400f0113
23e40173
402f0634
600f640c
00b30006
b00c602f
0026a00f
08040c56
602c21c3
6c4b6c6c
0a3432e4
301c0116
311c0b84
6c0c0000
36640266
08048056
23d22364
0053000c
2006002c
32e4602b
20260214
080401c3
61c3f016
602c72c3
646b2c6c
68d243c3
23c37fe5
446e2364
433c640c
606c2a1d
a5d2ad4c
24c316c3
566437c3
0f5604c3
00000804
405c3016
442b1804
672c200c
60277f85
315c06b4
6c0c0724
48802fcb
53c3700c
0ab425e4
0d24205c
0044323c
21946007
0075323c
302c0333
23e431c3
205c0ab4
323c0d24
60070024
323c1494
01930035
15c3b04c
0db421e4
0d24205c
0014323c
32c368f2
305c6072
606c0d27
36646c8c
08040c56
405c7016
c00c1804
205cbb2c
323c0d24
60070014
242b2d54
ffc0353c
06b46027
0724365c
afcb6c0c
708c2680
15e453c3
7f060435
01732383
0024323c
18546007
35c3b06c
061413e4
2583bf26
0d27205c
323c0193
6cd20044
53c3700c
083515e4
629232c3
0d27305c
6c8c606c
0e563664
00000804
ae243016
806cf524
4664902c
4004353c
f32462d2
08040c56
600c7016
0361335c
66d263c3
2fc30416
62c34385
ae242056
606cf524
36c38c2c
353c4664
62d24004
0e56f324
00000804
50c33016
506b846c
23e4704b
01160b94
0b84301c
0000311c
001c6c0c
366400a7
706b8056
523c500c
506b3b9d
602532c3
0c56706e
00000804
0136f016
041670c3
43052fc3
205682c3
235c600c
42d20361
515c244f
353c0293
c580180c
bfe5abd2
8d0c7c6c
163c07c3
4026fc4f
466438c3
8076fed3
08040f56
326431c3
6027402c
680c0394
63f200b3
0053682c
0c2b684c
00000804
600c3016
2d2c6c2c
533c68a0
6e32488c
205c6212
8d0026a4
253c300c
602601f4
200d233c
328331c3
505c65d2
100426f6
12a30073
0c56300f
00000804
600c3016
2d2c6c2c
533c68a0
6e32488c
205c6212
8d0026a4
253c300c
602601f4
200d233c
328331c3
32e365d2
700f3183
505c0093
100426f6
08040c56
3f36f016
91c360c3
c3c382c3
a05c802c
601004a4
0006b050
08cc78bc
fe00101c
28c39183
b00c43d2
b02c0053
ed6c786c
06c3e6d2
29c318c3
76643cc3
740b542b
199423e4
45d228c3
801cb02c
00930000
801cb00c
542b0001
23e4740b
786c0c94
09c36c6c
366414c3
282b2dc3
602531c3
0793682e
6c6c786c
14c309c3
542b3664
602532c3
236423c3
38c3542e
10946007
672c1bc3
25946087
215c64ac
8c6c0704
0b00301c
296b0c0c
46642d32
1ac30353
6007640c
065c1b54
60cc1804
21e413c3
60060535
680f2ac3
1ac30153
6ed2642c
13c360ac
0a3521e4
2ac36006
00d3682f
6c2c78ac
15c306c3
00063664
08cc82bc
0f56fc76
00000804
0336f016
81c350c3
802c92c3
04a4705c
0006d04c
08cc78bc
64d2782b
782e7fe5
08c307b3
300c0fd2
8007842b
01161a94
0b84301c
0000311c
02a66c0c
80563664
302c01d3
8df2842b
301c0116
311c0b84
6c0c0000
009d001c
80563664
057304c3
32c3442b
23c37fe5
442e2364
600738c3
74ac1e94
05c36c0c
02133664
1804355c
10c30cac
04b421e4
5c2f4026
0ccc00d3
21e410c3
402603b4
746c5c0f
05c36c4c
29c318c3
40c33664
00b30006
60077c2c
fe93e654
08cc82bc
c07604c3
08040f56
72c3f016
436440c3
04e4615c
1384515c
341c34c3
6ad24000
301c0116
311c0b84
6c0c0000
36640906
81c78056
812710b4
355c37b4
331c0a24
2a540200
00c7373c
6c4b7980
60476c32
05532394
fdc0343c
331c3364
12b40081
008c431c
431c0854
05b40094
088b343c
12946007
0095431c
431c0f54
1494009d
01160173
0b84301c
0000311c
08e66c0c
80563664
343c0133
03c30020
60860364
0a4d355c
343c0113
03c3ffe0
40460364
0a4d255c
08040f56
42c3f016
636460c3
736471c3
6dec696c
366402c3
045c50c3
340017a4
4010301c
0126640e
301c042e
644e0100
633c31c3
e4ae046e
06c3cc0b
1479645c
702c263c
345c4c0e
68121471
722c64ee
04c36c8c
366415c3
08040f56
80263016
40090213
033c30c3
3fc5009e
0bb401e4
035444a7
02944507
24208006
0c006025
f0b42027
0c5604c3
00000804
52c3f016
436440c3
636461c3
6dec696c
366402c3
155c70c3
008017a4
335c76ac
6e7204c3
62a6600e
740c602e
0624335c
606e6ee9
363c86f2
7fe50286
00f37f32
0286363c
7f3233c4
69a04066
8086608e
20c380ae
123c2206
30c3076e
043e433c
455c04c3
143c1479
2c0e702c
10c3080b
1471055c
40ac303c
762c680e
05c36c8c
366417c3
08040f56
0736f016
a0c3ff96
403781c3
e25743c3
90c34264
bfff941c
333c6297
275c00c7
ad0004e4
6dec7d6c
366407c3
375c60c3
018017a4
335c7eac
6e7204c3
20c6600e
343c202e
604e400c
323c4017
606e442c
602620c3
056e323c
34c394c9
0018341c
04946107
0101101c
20c3280e
046e923c
620610c3
076e313c
335c7c0c
303c03e1
880b066e
475c54c3
343c1479
680e72ac
25c3a40b
1471575c
412c353c
393c640e
3364f480
05356187
341c3ac3
64d24000
6872600b
7e2c600e
07c36c8c
366416c3
e0760196
08040f56
0f36f016
b0c3fd96
43c362c3
525c2970
57cb1384
0060323c
359d753c
355c29d2
331c0a24
04940200
0010323c
37c377ce
60073164
355c0f15
647209c3
09c6355c
7fff741c
0053a55c
0000801c
60b76026
a55c00f3
801c0043
20060001
798c20b7
341c6c0c
65d20008
0000801c
40b74026
60073bc3
19c31154
07c3652c
366416c3
8077c037
880c29c3
212607c3
7f5c2ac3
37c30041
18c34664
11542007
894c29c3
20260bc3
36c34006
74e94664
79c368d2
00069d4c
40262006
466436c3
f0760396
08040f56
fe967016
d56ca00c
09a3355c
155c2006
612709a6
61470454
06d35694
04e4355c
2c29592c
2d0941c3
722c013c
266415c3
04e4355c
42c34c29
323c4d09
a037722c
80778006
03c3980c
21c32146
46646026
1384355c
0100101c
0a27135c
1384255c
09c3425c
341c34c3
325cffcf
255c09c6
325c1384
687209c3
09c6325c
05c3798c
36643fe6
358c0413
323c440c
65d20084
639232c3
0093640f
05c3788c
355c3664
602713a1
75cc0694
05c36c2c
00d33664
6c4c75ac
15c30006
355c3664
48061384
0a27235c
0e560296
00000804
405c1016
41e61384
0ab6205c
6e8c606c
245c3664
32c309c3
feff341c
09c6345c
08040856
1384205c
09c3125c
341c31c3
00060003
11946067
0a24225c
2006323c
0b0d333c
fff0133c
4006323c
0b0d333c
31a37fe5
f88c033c
00000804
41c37016
c56c0364
1471215c
17c7323c
0564215c
6e8c6d00
a2864c2c
66d2684b
48e979cc
03643664
700ca506
0d89235c
20c349d2
4000241c
16944007
14b401c7
345c00f3
61c709e4
01c70635
790c04b4
00f302c3
08b461c7
063501c7
0026790c
24c315c3
0e563664
00000804
0336f016
50c3ff96
905ce16c
648c0584
0079835c
1384405c
305c6006
648c13a5
788bc980
0976345c
33647fe5
0a356ee7
4006606c
8dec4037
4e262386
46646006
36c30813
053f233c
0a06245c
03e0043c
245c13c3
b0bc0973
600608cb
09f6345c
32c35849
0010341c
12546007
09c3245c
341c32c3
66f20002
0a24345c
0004341c
7d6c64d2
366405c3
345c6026
383c09f6
333c208c
29c30cc7
68d269a2
06546047
32c35849
0001341c
60266cd2
13a5355c
09f3245c
345c46d2
607209c3
09c6345c
01960006
0f56c076
00000804
fe96f016
e16c50c3
1384405c
c980648c
335c62ac
04c30524
233c16c3
b0bc0300
245c08cb
32c309c3
0002341c
7d6c64d2
366405c3
64d2782b
00ff341c
301c0073
345c00ff
50c909e6
7fe532c3
3f5c6077
62e70021
746c0b35
40374006
05c38dec
4de62386
46646006
345c03d3
584b09c3
607245d2
09c6345c
609200f3
09c6345c
05c37d6c
60063664
400673ce
09a7245c
09c3245c
341c32c3
345cfffb
600609c6
09f6345c
02960006
08040f56
3f36f016
b0c3fe96
126453c3
d2c32037
935cd264
135c1384
313c1471
c3c317c7
0564255c
4cc3c284
6c2c728c
756c6077
05c36dec
a0c33664
680c558c
0004341c
682c67d2
01f1835c
03f0733c
09c300d3
0973805c
03e0793c
1ac376ac
04c4235c
455c6500
ce0017a4
00070bc3
9d8b1494
11548007
06c38832
430617c3
08cbb0bc
00c6b65c
01a0343c
c345fd80
283c84a4
0053fe60
06c328c3
b0bc17c3
1dc308cb
063c28d2
1c3c0040
40c60480
08cbb0bc
236428c3
435c76ac
6a0004c4
638e0ac3
135c76ac
688004c4
401760ce
608645d2
8000311c
4ac3620f
17a4055c
558c3000
341c680c
60070004
682c1354
01f1335c
640e6e72
0600201c
301c444e
646e0205
6c2c758c
40066c2b
1d356207
49c30313
0973345c
640e6e72
1800001c
201c044e
446e0205
0a03245c
5804323c
13cb6cf2
60a530c3
359d343c
053561c7
008b001c
0053048e
4057448e
45d2484b
345c49c3
64ae0a49
033c31c3
40c3043e
1479055c
722c203c
355c4c0e
68121471
762c64ee
05c36c8c
36641ac3
680c558c
680f6292
fc760296
08040f56
ff96f016
51c360c3
415ce56c
045c1384
30c309c3
0003341c
84dc6067
345c0008
60870a24
000832dc
05546807
331c0026
7d940100
301c0006
311c0fe4
2cac0000
0873b4bc
32c353cb
343c60c5
6007351d
30ab0515
0a16145c
508b0093
0a16245c
70c953cb
051423e4
05c37d6c
0bd33664
0a13145c
508c263c
00a0313c
13b423e4
1323355c
08546027
12e4055c
028d333c
31e46a32
345c0434
65d20bd9
09f3645c
1854c007
045c0026
7c8c0bdd
366405c3
05c37d8c
111c22c6
3664000a
0200101c
0a27145c
155c0266
00bc1341
00260873
558c05d3
433c680c
80070084
682c2254
0981235c
002502c3
1f5c0037
135c0001
758c0985
325c4c2c
60a70981
7c6c05b4
366405c3
325c0193
65720993
0996325c
335c746c
140c0824
366416c3
00f306c3
05c37c6c
04c33664
00060053
0f560196
00000804
40c37016
1384205c
a06cc16c
125c2006
305c0bdd
135c1384
31c309c3
0001341c
60a662d2
09c6325c
125c2086
40060a27
0ab6245c
04c3768c
75ac3664
21e604c3
345c3664
20061384
0bd5135c
6c2c71ac
366404c3
145c0266
b8bc1341
02660872
1341145c
087300bc
04c3798c
36643fe6
08040e56
0136f016
50c3ff96
1384405c
0170e06c
145c2006
305c0bdd
235c1384
32c309c3
0001341c
13546007
345c6026
53cb09c6
23e470c9
345c0554
61070a24
758c0c94
341c6c0c
c0260008
00b367d2
09c6345c
005363c3
345cc006
61070a24
355c0a94
235c1384
32c309c3
0001341c
3c946007
73ce6006
145c2006
355c0a27
602713a1
345c0b94
68d209f3
09c3145c
341c31c3
345cfffe
400609c6
09f6245c
301c0006
311c0fe4
2cac0000
0873b4bc
155c0266
00bc1341
60060873
0ab6355c
05c37e8c
7dac3664
21e605c3
355c3664
20061384
0bd5135c
6c2c75ac
366405c3
698c28c3
3fe605c3
746c3664
142c6dcc
40862026
30c33664
6bf23264
6106cad2
0a27345c
155c0266
2cbc1341
01f30873
155c0266
b8bc1341
c9d20872
20372006
05c39dec
42e62026
46646006
80760196
08040f56
0736f016
a00c90c3
946cf56c
655c1430
055c1384
05f21469
13a1355c
54946027
0a24365c
0200331c
331c0754
42541000
54946107
5bcb09f3
23e478c9
01160a14
0b84301c
0000311c
09466c0c
80563664
08c371cc
40862006
30c33664
60073264
51d01554
1804255c
045c49c3
30c30361
7f327fe5
080c933c
202608c3
894b39c3
a6644e00
326430c3
7c6c63f2
9dac0493
10c30026
600625c3
02664664
1341155c
0872d0bc
8000001c
0000011c
0a27065c
101c0353
165c2000
9d4c0a27
20060006
35c34026
02664664
1341155c
0872b8bc
7d6c0153
366405c3
026600d3
1341155c
0872d0bc
0f56e076
00000804
50c33016
6ccc606c
2006000c
40c33664
335c76ac
255c04c4
2d0017a4
08cb9cbc
235c76ac
538e04c3
17a4255c
708f7100
235c76ac
50ce04c3
70ee6006
70af6006
245c4086
718f01d5
1471355c
01ed345c
1479255c
027d245c
0c5604c3
00000804
0336f016
505c40c3
005c1384
145c0564
255c1471
323c09c3
60070024
355c7894
341c0a24
60071000
323c7294
60070014
313c6e54
c18017c7
341c780c
64d20001
1469245c
345c45f2
602713a1
8ebc6094
70c30895
0bb3065c
09a4355c
755c64f2
0ab309a7
83a487c3
93c3744b
4240301c
000f311c
328d693c
0bb486e4
09d3155c
09e3255c
03e46880
68000434
04b431e4
03e4740b
355c0eb4
60870a24
355c0a54
67f209f3
13a1345c
31946027
2f3586e4
09d6055c
0a24355c
03546087
09a7755c
145c0266
a2bc1341
41e60872
0ab6245c
6e8c706c
366404c3
13a1345c
03946027
00f371cc
1384345c
235c4026
71ac0bd5
04c36c2c
355c3664
617209c3
f7fb201c
355c3283
680609c6
0a27355c
0f56c076
00000804
0336f016
50c3fc96
92c361c3
e2d783c3
628c0357
600743c3
6c091454
400660f7
04946027
00613f5c
00d723c3
361c30c3
7fe50003
02c37f32
00b703a3
00414f5c
163c05c3
265c0d40
34c30784
091498bc
240b2317
0696165c
00c0201c
46c3582e
17c4355c
1f866065
380b3083
76ac45a0
0404335c
30836065
343c4980
323c604e
700f601b
17c4355c
30836065
765c83a4
29c306e7
3a544007
365c60a6
700c0286
323c40a6
700f231b
104d0066
200637c3
0040111c
60073183
973c1a54
373c03f4
60070034
56ac1454
0404325c
1f866065
125c3083
6c8004c4
71803884
0020033c
29c313c3
090a5abc
00534046
76ac4006
0404335c
1f866065
18c33083
6d006580
2f5c6077
508d0021
60860533
0286365c
4086700c
231b323c
0046700f
76ac104d
0404335c
3f866065
83843183
00078f5c
00013f5c
055c708d
11ed09e1
17c4355c
31836065
59806185
335c746c
05c30764
482b280b
065c3664
255c0686
265c09e1
355c0705
000617c4
0060011c
20c37083
139472e4
1f866065
61853083
746c5980
0764335c
280b05c3
3664482b
065c0364
055c0686
00932947
165c2006
57660686
070d265c
c0760496
08040f56
0336f016
50c3ff96
82c391c3
e06c8364
c037c506
21669fcc
32c34006
40c34664
355c56ac
606517c4
31833f86
04a4125c
01806c80
188419c3
b0bc26c3
375c08cb
05c30404
366414c3
c0760196
08040f56
40c31016
0724105c
19542007
0704345c
100462f2
345c7fe5
345c0707
6c2c0724
0727345c
345c63f2
706c0747
05a4335c
366404c3
0724145c
e9942007
08040856
3f36f016
50c3fc96
82c391c3
60708030
21c3a250
111c2006
21830040
45544007
400609c3
0020211c
00070283
355c1b54
606517c4
31833f86
458018c3
65052a8b
636463c3
00a0363c
a8c328c3
6b00a384
32c34c4b
0001341c
e1068006
48946007
49c30313
311c6006
43830100
13548007
17c4355c
3f866065
18c33183
290b4580
63c36205
363c6364
a8c300a0
40c3a384
05d374c3
301c0116
311c0b84
6c0c0000
36640d66
04138056
600649c3
0200311c
80074383
305c1054
606517c4
31833f86
63c36185
363c6364
a8c30060
12c3a384
01b38026
301c0116
311c0b84
6c0c0000
36640d86
14c38056
a1c364c3
313c71c3
610700c4
80070454
0008d2dc
200639c3
0090111c
31e43183
355c7494
606517c4
32835f86
658018c3
233c6c2c
7f86708c
43f22383
0564255c
0564155c
76ac48a0
0444335c
3230141d
17c7333c
eed22580
67326409
155c6bf2
21c30949
40f74025
00613f5c
094d355c
640c0bb3
0002341c
155c6bf2
21c30951
40b74025
00413f5c
0955355c
155c09f3
21c30959
40774025
00213f5c
095d355c
1254e007
200639c3
1000111c
6cd23183
0961355c
08b46087
0010233c
3f5c4037
355c0001
1bc30965
0cc365cc
40c62026
30c33664
60073264
393c2954
2dc31e8b
05c3882c
27c32006
3ac323a3
e0074664
39c31d54
111c2006
31831000
16546007
255c4006
02530965
65cc1bc3
20260cc3
366440c6
326430c3
88f269d2
2dc3e7f2
05c3684c
26c318c3
04963664
0f56fc76
00000804
3f36f016
40c3f996
c2c3b1c3
04a4005c
300c00f7
2bc32177
6312682c
6c00080c
324ccc2c
345c21b7
606517c4
32835f86
6006f981
37c36137
011c0006
30837c00
345c64d2
6cd20a44
642c20d7
37c369f2
211c4006
32834000
f2dc6007
37c30009
011c0006
30834000
345c67d2
4c4c2544
4c4f4025
37c30213
111c2006
31832000
2544245c
682c65d2
682f6025
68ac0093
68af6025
682c40d7
13546007
2544245c
6025686c
0157686f
6087632c
305c0a94
40060724
0135235c
0724305c
0d4f0006
200637c3
1c00111c
6dd23183
400637c3
6000211c
67f23283
616c0197
17c304c3
366426c3
200637c3
0200111c
65d23183
694c4197
366404c3
000637c3
0360011c
60073083
20c31554
125432e4
011c0006
10c30120
0c5431e4
40066006
0340211c
00067283
0240011c
71e410c3
60260294
419765d2
04c3694c
0bc33664
6312602c
ac80200c
6007742a
01160a74
0b84001c
0000011c
0d06600c
80563664
642c1bc3
0010233c
345c442f
23e40941
40060394
345c442f
606517c4
30831f86
2006542c
201c2d61
540e0200
30c3142b
4000341c
6007342e
2e13d394
0116eaf2
0b84201c
0000211c
08a6680c
80563664
2544345c
40254c0c
37c34c0f
011c0006
30830360
16546007
32e420c3
00061354
0120011c
31e410c3
40060d54
000637c3
0340011c
20063083
0240111c
30e401c3
40260294
219745d2
04c3654c
d01c3664
a01c0001
9ac30000
2bc38ac3
6312682c
ac00080c
6007742a
01160a74
0b84201c
0000211c
0d26680c
80563664
0009a31c
72ac1254
0404335c
1f866065
101c3083
65a00fff
075493e4
602c00d7
38c383a3
36546007
682c40d7
01576ed2
6087632c
305c0a94
40060724
0135235c
0724305c
0d4f0006
17c4345c
3f866065
542c3183
0d610006
0200101c
542b340e
141c12c3
60064000
0bc3742e
233c602c
402f0010
0941345c
0000d01c
0001801c
7d9423e4
2bc36006
d3c3682f
0001801c
542c0ed3
00070ac3
584f1694
21c3340b
345c4185
606517c4
30831f86
78ce6980
21c3340b
345c4185
606517c4
92c33083
06539384
00103a3c
3f9d263c
0003855c
335c72ac
09c30404
00370884
0030133c
12835f86
0fff301c
60776ca0
180c0a3c
23c36017
23e46057
78000734
0066835c
9084140b
58000233
321c31c4
39a40fff
72ac68ce
0404335c
3f866065
201c3183
92c30fff
706c93a4
01576ccc
36642026
142f20c3
17c4345c
1f866065
20063083
201c29e1
540e0200
6006342b
0bc3742e
233c602c
402f0010
0941345c
049423e4
2bc36006
141c682f
2a3c4000
40b70010
00413f5c
a264a3c3
0000801c
04dc2007
a65cfff3
37c30296
011c0006
30830200
3e546007
0006965c
20071dc3
345c5354
60250704
0707345c
0744345c
645c64f2
00530727
645ccc2f
40060747
37c3582f
011c0006
30830080
42546007
642c1cc3
0724245c
644c63d2
3cc30053
145c4c2f
0cc30744
600c204f
0704245c
600f6d00
345c6006
345c0727
345c0747
245c0707
682c25a4
682f6025
01370026
965c0433
1dc30006
16542007
680c2cc3
680f6025
63f2684c
0053c82f
3cc3cc2f
0006cc4f
345c182f
4c2c25a4
4c2f4025
21372026
706c00f3
05a4335c
16c304c3
2bc33664
6312682c
6c00080c
6c2a2c2c
10156007
345c61c3
606517c4
30831f86
37c3e581
111c2006
3183c000
a4dc6007
4117ffdc
008646d2
1341145c
0872a2bc
211c4a86
60262010
6f86680f
2010311c
0c0f0026
2c0f2086
2bc3280f
6312682c
6c00080c
6c2a2c2c
32e44006
345c0715
606517c4
32835f86
32c34581
011c0006
3083c000
004666f2
1341145c
0872b8bc
fc760796
08040f56
311c6f86
40462010
201c4c0f
211c817e
680b2010
dfff341c
680b680e
bfff341c
201c680e
211c817c
680b2010
dfff341c
680b680e
bfff341c
301c680e
311c806a
201c2010
4c0e00e0
305c6026
0804051d
311c6d06
40462010
201c4c0f
211c817e
680b2010
6d723364
680b680e
6e723364
201c680e
211c817c
680b2010
6d723364
680b680e
6e723364
301c680e
311c806a
201c2010
4c0e0160
305c6006
0804051d
0736f016
2006fd96
c00c20b7
0684765c
5c095870
1094101c
0020111c
933c6880
323c400c
133cfff0
2077f88c
00212f5c
19c35c0d
201c644b
211cffff
12c30000
495431e4
0104201c
3ac34037
06c38fcc
400621c6
466432c3
365c80c3
606517c4
31833f86
74eba180
74ee6072
0104201c
365c544e
606517c4
62053183
8ebc8180
34c30895
027f033c
19c303c3
0100201c
08cbb0bc
47d25c2b
ffaa301c
0000311c
00d360b7
ffbb101c
0000111c
053c20b7
1f3c0060
40860080
08cbb0bc
325c580c
60250544
0547325c
325c2ac3
06c30404
366418c3
165c00c6
b8bc1341
7c2b0872
20066dd2
40063c0d
301c5c2e
311c8180
101c2010
2c0e4000
301c0113
311c8180
201c2010
4c0e2000
817e201c
2010211c
341c680b
680e9fff
e0760396
08040f56
0f36f016
70c3fd96
52c3a1c3
9f5c0397
8f5c0183
400601a1
d40b5c0d
400640c3
133c40b7
3f5c0804
60370041
0fc3345c
239436e4
0fd3245c
23e4742b
245c1e94
744b0fe3
199423e4
345c28d2
331c0ff1
135400ff
119438e4
323c4097
61800147
1003335c
40774026
0f9439e4
00212f5c
60065c0d
01336077
32c34097
60b76025
60678285
0473d194
b3c36017
0002b31c
3f5c1eb4
2ac30001
4017680d
0147323c
543c8180
340c2040
60076057
606c1054
05a4335c
40063664
6006540f
1006345c
245c5fe6
7fe60ff5
0fc6345c
f0760396
08040f56
50c37016
603c40c3
145c03c0
20071024
746c1154
05a4335c
366405c3
345c6006
345c1027
7fe61006
0ff5345c
345c7fe6
82850fc6
ea9446e4
08040e56
6ca06406
318d003c
00000804
118d003c
00000804
20c330c3
ff00101c
ff00111c
48322183
00ff101c
00ff111c
033c3183
0804412c
3f36f016
00b7fb96
607702c3
636461c3
815c2097
21c30013
42c32884
0f4f343c
433ca4c3
80f7fff4
800c72c3
173ca02c
4103084e
222604c3
08f506bc
96005003
10bc04c3
500308f5
04c39600
06bc2066
500308f5
04c39600
0cbc2046
500308f5
5c2c9600
04c34203
06bc2226
500308f5
04c39280
08f510bc
92805003
206604c3
08f506bc
92805003
204604c3
08f50cbc
92805003
43037c4c
222604c3
08f506bc
92805003
10bc04c3
500308f5
04c39280
06bc2066
500308f5
04c39280
0cbc2046
500308f5
363c9280
430300f4
222604c3
08f506bc
92805003
10bc04c3
500308f5
04c39280
06bc2066
500308f5
04c39280
0cbc2046
500308f5
101c9280
111caaaa
41030003
222604c3
08f506bc
92805003
10bc04c3
500308f5
04c39280
06bc2066
500308f5
04c39280
0cbc2046
65c308f5
53006003
533c7c6c
05c3811c
06bc2226
46c308f5
b6004003
10bc05c3
400308f5
05c3b600
06bc2066
400308f5
05c3b600
0cbc2046
400308f5
4097b600
31c328cb
38a47c45
736473c3
32c340d7
83c37e45
60068164
63c3c3c3
11936137
0034973c
108cb73c
e006dac3
2dc30433
0004d21c
5303680c
222605c3
08f506bc
b2804003
10bc05c3
400308f5
05c3b280
06bc2066
400308f5
05c3b280
0cbc2046
400308f5
373cb280
73c30010
7be47364
38c3df14
2b3c39a4
6d00130c
d364d3c3
81648dc3
0000831c
01160c15
0b84201c
0000211c
001c680c
36640089
00b38056
63f238c3
09933bc3
25d219c3
3ac32bc3
299d633c
00102c3c
3f5c4037
c3c30001
3c3cc264
20970010
3e1da13c
180c3c3c
eccb6580
400729c3
1ac32e54
633c640c
e027832c
602604b4
04b36137
150316c3
01c351c3
06bc2226
400308f5
05c3b600
08f510bc
b6004003
206605c3
08f506bc
b6004003
204605c3
08f50cbc
b6004003
0002a21c
ffe0373c
736473c3
ffe03d3c
816483c3
18c33bc3
34dc2007
4117fff7
1ac344f2
3a1d613c
32c340d7
341c60c5
60270003
66d20a54
0d546047
1c946067
561c0233
0313005a
0ff4363c
5a00351c
02535303
ffff641c
211c4006
62a3005a
301c0153
311cffff
638300ff
111c2006
61a35a00
05c35603
06bc2226
400308f5
05c3b600
08f510bc
b6004003
206605c3
08f506bc
b6004003
204605c3
08f50cbc
b6004003
222605c3
08f506bc
b6004003
10bc05c3
400308f5
05c3b600
06bc2066
400308f5
05c3b600
0cbc2046
24c308f5
75002003
700f8057
0596502f
0f56fc76
00000804
3f36f016
60c3ea96
73c3b1c3
0f5c0006
0f5c02bd
200602b5
24b72477
17c4335c
0030233c
7f8612c3
78801383
533c6c2c
1f86708c
a3b75083
533c740c
a177288b
01b70706
03156007
a1b7a306
04371c6c
0320313c
a384a6c3
23837f86
925c5900
abeb0143
0804393c
00ff001c
637702f7
225c67d2
43770203
000f241c
400642f7
02a6265c
62776006
00f4353c
802663f2
393c8277
00064004
66f202b7
165c2086
402602a6
625742b7
62dc6007
82970009
24dc8007
00860009
02a6065c
1003175c
275c2bd2
48d210a3
1143375c
80a665d2
02a6465c
7d4c6073
00065f5c
01610f5c
00250f5c
8c0ce0b7
05600f3c
05701f3c
39c32ac3
375c4664
61f71003
175c6ad2
31c310a3
233c7fe5
6046f88c
61f76d20
00e12f5c
02bd2f5c
343c81d7
7d800147
1027635c
02b90f5c
0147303c
353c5d80
325c0010
1f5c1006
313c02b9
7d800147
01612f5c
0ff5235c
02b94f5c
0147343c
5ac37d80
535cb40b
0f5c0fc6
303c02b9
7d800147
242b1ac3
0fd6135c
02b92f5c
0147323c
4ac37d80
435c904b
275c0fe6
3f5c0f81
48d202b9
0147333c
a0067d80
1056535c
333c0133
7d800147
1056235c
075c0c86
180b0f96
02b93f5c
0200031c
333c0894
7d800147
235c4006
51d31046
0147333c
203c3d80
301c1ff4
6d200200
1046315c
801c5073
8f5c0000
625701e7
14dc6007
7d4c0020
00065f5c
01614f5c
00254f5c
8c0ce0b7
05600f3c
05701f3c
39c32ac3
5f5c4664
a5f202b1
065c0026
4c9302a6
02b91f5c
0147313c
425c5d80
34c31003
325c6025
5f5c1006
353c02b9
7d800147
1024835c
03f43b3c
0020133c
17c4375c
1f866065
233c3083
313c0280
698007c4
d364d3c3
32c3580b
c3c33da4
a297c364
c2dca007
09c3000f
341c30c3
60074000
000f52dc
31c32157
000a341c
e2dc6007
3bc3000e
211c4006
32830001
64dc6007
c31c000e
67b40008
4cc36106
15c3ae20
08c31364
60a0000b
680e28c3
0980682b
233c600c
48a0600b
601b323c
9f3c600f
48c30440
0293045c
7fe530c3
71806312
53e46ccb
01162735
0b84301c
0000311c
08c66c0c
80563664
0293245c
fff0123c
180c313c
0ccb7180
323c9420
6312ffe0
698028c3
063e233c
003c08c3
28001e1d
4c0e4a20
19c30620
b0bc24c3
b62008cb
28c39484
0293125c
fff0313c
69806312
063e233c
443c48c3
2a001e1d
4c0e4aa0
19c306a0
b0bc25c3
78cb08cb
6c00184c
0ca01cc3
2a8029c3
b0bc2cc3
602608cb
28b363f7
ff803c3c
c364c3c3
0293265c
4b354027
fff0323c
39806312
063e913c
0007931c
49c31035
2e1d563c
035c7280
0477ffc4
ffe4235c
840b44b7
7f0534c3
07f3640e
59c36106
323c8ea0
6312ffe0
033c7980
4220063e
165c4c0e
313c0293
5f3cffe0
63120440
4ccb7980
05c33fe5
1e1d363c
24c32980
08cbb0bc
a484a5c3
0293165c
7fe531c3
79806312
063e433c
29a424c3
365c4c0e
0ac30293
3e1d163c
b0bc29c3
01f308cb
b84c58cb
035c6a80
0477ffc4
ffe4135c
323c24b7
78ceff80
0124af5c
0293265c
fff0323c
79806312
83f78026
a007accb
04171594
07c360ec
2e1d163c
36644026
0293165c
7fe531c3
0296365c
43f74026
a01c00b3
af5c0000
5cc301e7
900b48c3
58c37600
142b740e
640c3400
600b233c
51004cc3
601b323c
5f5c640f
353c02b9
7d800147
1043935c
105c08c3
21c30291
41375fe5
00813f5c
b264b3c3
34c398cb
53c33da4
49c35364
2d3c1293
323c424b
363c0010
62373e1d
323ca5f2
7980180c
8007accb
b31c2e94
0b940005
101c0116
111c0b84
640c0000
008a001c
80563664
68cc4417
20261c0c
20c33664
00104b3c
0f5c80f7
b0c30061
3b3cb264
18c30010
3f9d213c
180c3b3c
80066580
a2c38cce
0293015c
602530c3
0296315c
0200401c
180c3b3c
073554e4
698028c3
063e033c
00d35000
658018c3
063e033c
4c0e5400
2bd219c3
00103b3c
323c28c3
321c3e1d
a3c30200
00b3a9a4
0200101c
a3846620
103554e4
62200cc3
c364c3c3
71002dc3
63373364
762024c3
536453c3
94c38006
25c303f3
62a00cc3
c364c3c3
74000dc3
63373364
43c372a0
1cc34364
0f5c28f2
303c02b9
7d800147
1046435c
23f219c3
00d359c3
62a009c3
936493c3
1d3ca006
0ac31ff4
25806217
08cbb0bc
0184df5c
00070cc3
fff6b4dc
20072297
42577954
71944007
02a3465c
341c34c3
365cfffb
a3d702a6
4054a007
30c30397
24176105
07e4415c
435708c3
a19712c3
3f3c4e80
466404c0
04d76457
31e410c3
64970694
42c34517
285434e4
355ca417
07c305a4
366418c3
02b90f5c
0147303c
20067d80
1027135c
02b92f5c
0147323c
80067d80
1006435c
02b95f5c
0147353c
1fe67d80
0ff5035c
02b91f5c
0147313c
5fe67d80
0fc6235c
4f5c05b3
343c02b9
7d800147
535ca006
0f5c1027
303c02b9
7d800147
135c2006
2f5c1006
323c02b9
7d800147
435c9fe6
5f5c0ff5
353c02b9
7d800147
035c1fe6
24170fc6
0404315c
18c307c3
00d33664
02a3365c
365c6172
169602a6
0f56fc76
00000804
311c6a86
20862010
205c2c0f
40070a61
40061454
0504305c
0200101c
2f1d133c
180c323c
0504105c
20066c80
40252c2e
0941305c
ef1423e4
00000804
0336f016
301cfe96
311c0bb4
8c0c0000
06a4845c
0664745c
611cca86
580c2010
311c6f86
ac0c2010
780c5283
0010341c
712c67d2
04c36cec
22063664
35c3380f
211c4006
32830010
1b546007
2524245c
6025692c
345c692f
2ce904c4
341c31c3
66d20001
6ccc712c
366404c3
01160153
0b84301c
0000311c
0e066c0c
80563664
0024353c
712c65d2
04c36c2c
353c3664
6ad20014
0484345c
345c6025
712c0487
04c36c4c
35c33664
ff00201c
000f211c
60073283
345c1154
60250464
0467345c
2524245c
6025682c
712c682f
04c36c6c
25c318c3
353c3664
6ad20044
2524245c
6025686c
712c686f
04c36c8c
353c3664
60070084
201c1054
211c0448
680c2010
680f6092
311c6a86
21062010
680c2c0f
680f6072
0404353c
23546007
dcbc04c3
245c0910
688c2524
688f6025
1471245c
17c7323c
0564145c
6c0c6c80
0001341c
245c6bd2
48d21469
13c37f89
20772025
00212f5c
6a865f8d
2010311c
2c0f2806
0804353c
712c66d2
04c36cac
366418c3
0204353c
34546007
2524245c
602568cc
201c68cf
211c0090
680c2010
fff4633c
501c0006
511c7300
e0262010
173c92c3
31c3000d
60073683
29c31754
303c280f
145c03c7
6c8006a4
315c2d0c
69d201f9
fff0833c
00078f5c
00012f5c
01fd215c
3364740b
0025740e
0187a085
201ce194
211c0090
680c2010
2000341c
13546007
2000101c
245c280f
68ec2524
68ef6025
301c0116
311c0b84
6c0c0000
008f001c
80563664
c0760296
08040f56
0736f016
60c3fa96
0070a1c3
1504705c
06c4905c
1469005c
46540007
1471165c
17c7313c
0564265c
6c0c6d00
0001341c
3a546007
0c73065c
341c30c3
60070010
8ebc3354
20c30895
15c4165c
065c6080
2c2015a4
15c7165c
15a7265c
1583365c
12e4265c
228d333c
1e3513e4
335c780c
341c0504
6dd20001
165c2206
786c1666
40374206
06c38e0c
00c5101c
46646006
60376006
81ec08c3
218606c3
466423c3
165c2006
5d0915c7
6d544007
09e4365c
69546007
60077d29
79cc2c94
06c36c0c
2a123c2b
36644026
465c50c3
1c2b1771
5cbc14c3
303c0a7c
141d500c
133c3530
343c0010
1383fff0
3f5c20f7
61370061
00810f5c
3d491c2d
265c2c80
32c31771
13837fe5
1f5c20b7
3c2d0041
5d2d4026
303c1c29
165c0cc7
6c800584
0641235c
1c544007
0604365c
44724c6c
1c2c4c6f
2c6c39c3
301c4046
311c0fe4
6cac0000
08745abc
005c0ac3
0df21503
315c18c3
06c30744
36643c29
365c00d3
4d0c2524
4d0f4025
32c35c29
60776025
00210f5c
1f5c0177
3c2d00a1
1771365c
03d430e4
7c2d6006
305c08c3
06c30504
6a863664
2010311c
0080101c
06962c0f
0f56e076
00000804
0f36f016
90c3ff96
72c381c3
ff00301c
000f311c
673c7383
b01c408c
b11c0b84
a01c0000
04d30001
0cbc06c3
50c308ce
03c7303c
898028c3
602770cb
01160854
680c2bc3
00a0001c
80563664
500d3a3c
638333e3
23c37029
00fd241c
3f5c4037
702d0001
0070053c
125c29c3
00bc1341
c0070873
6d06da94
2010311c
0196ec0f
0f56f076
00000804
305c10c3
4c0c2524
4c0f4025
0a61005c
00460cf2
1341115c
0872a2bc
311c6d06
40262010
03334c0f
311c6a86
00262010
40060c0f
0504315c
0200001c
2f1d033c
180c323c
0504015c
00066c00
40250c2e
0941315c
ef1423e4
00000804
301c10c3
311c8182
6c0b2010
236423c3
341c32c3
60076000
32c31754
4000341c
305c65d2
40260684
201c4c2e
211c817e
680b2010
351c3364
680e6000
115c00c6
a2bc1341
08040872
40c31016
301c01c3
311c08cc
2c0c2010
6c0c6085
706c47d2
0524335c
366414c3
200f0073
0856602f
00000804
ff963016
6037640c
6e20880c
40c3600f
282c642c
543caca0
4017027e
600c2006
023532e4
74a02026
0196700f
08040c56
ff963016
12c341c3
4037500c
6d00640c
50c3600f
502c642c
453c8d00
4017027e
600c2006
023432e4
70802026
0196740f
08040c56
1364ff96
3f5c2037
305c0001
0196016d
00000804
4c6c600c
06a4225c
0544035c
26642026
00000804
0066600c
1341135c
0872a2bc
00000804
1341305c
13c30066
087300bc
00000804
335c600c
201c1341
211c0fe4
27d20000
13c30026
d4bc490c
00d308c8
13c30026
b8bc490c
080408c8
0136f016
50c3fe96
605c72c3
848c06a4
0ad211e9
301c0116
311c0b84
6c0c0000
36640b86
51e98056
141c12c3
313c000f
055c00c7
6c0004e4
4c0d4026
0c2d1109
4c4d5129
80c31149
203c1169
4c4e442c
4ccd51c9
20c311e9
000f241c
0f5c4077
0ced0021
483250cb
0f5c4037
0d0d0001
36c35380
880b0006
882b8c4e
884b8c6e
886b8cae
00258c8e
67854105
f4940187
335c746c
05c306e4
00263664
80760296
08040f56
1f36f016
60c3ff96
82c3c1c3
407093c3
40076010
323c3054
533c080c
a037928d
87cc1ac3
40862026
46646006
365c70c3
531c17c4
093500ff
3f866065
61803183
40724ceb
ac4e4cee
4ccc780c
17c4365c
3f866065
62053183
60377d80
0bc3882c
28c31cc3
466439c3
325c2ac3
06c30404
366417c3
f8760196
08040f56
0336f016
e00c62c3
945c848c
50eb0049
341c32c3
833c000f
341c0034
64d20001
6dcc60cc
53003664
01532006
0006680c
4130011c
082c6c00
41450c0f
19e42025
383cf614
65d20024
6c6c7ccc
366407c3
c0760026
08040f56
1f36f016
60c3ff96
607092c3
e48c4010
875c9d09
3ceb0049
341c31c3
c33c000f
341c0034
64d20001
6dcc60cc
343c3664
533c828d
a037080c
8bcc2bc3
202606c3
60064086
40c34664
17c4365c
00ff531c
60650935
32835f86
4ceb6180
4cee4072
39c3ac4e
365c5d80
606517c4
3583bf86
31806205
01f30006
a006680c
4130511c
ac0c6e80
680ba42f
a82b640e
4145a42e
00252145
f11408e4
00243c3c
5ac366d2
6c6c74cc
36640ac3
315c1bc3
06c30404
366414c3
01960006
0f56f876
00000804
00000804
335c606c
36640424
08040006
f0963016
0fc350c3
8024101c
0012111c
e6bc4806
4fc308cb
32c3500c
039453e4
01130026
2f3c8085
32c30400
f59443e4
10960006
08040c56
13643016
536452c3
60ec800c
245c26d2
46f20519
00536c4c
04c36c2c
a0073664
345c1754
60070519
301c1354
311c8180
201c2010
4c0e4000
2000201c
201c4c0e
211c817e
680b2010
9fff341c
0c56680e
00000804
ff96f016
01c360c3
65e9248c
17c7533c
0564365c
84eb6e80
141c14c3
2037000f
00017f5c
02ad735c
4880208c
0564365c
60262e80
0406315c
415c880b
32c30416
013e733c
0426715c
015c0c0b
8c0b04b6
0486415c
715cec0b
084b0496
0436015c
343c42c3
6132033e
03c37fe5
315c0364
30e40443
60060454
0466315c
0446015c
715ce88b
08ab04e6
0506015c
315c68cb
41c50456
01d32006
0520313c
765c6112
6f800564
159d023c
313c0ec1
13c30010
700b1364
f1b431e4
01960006
08040f56
0f36f016
0584505c
6509248c
652943c3
422c233c
0024823c
0100713c
0806323c
09cbb33c
6bc385e9
c5c9cdd2
17c7363c
105c93c3
91840564
0cc7343c
49c31580
343c00f3
15800cc7
0b80403c
323c9bc3
a1460204
0000a01c
22946007
0104323c
6007a026
323c1d94
64d20084
a086e025
323c00d3
66d20044
5ac3e025
0001a01c
123c01f3
a2060404
700c2bf2
44f228c3
085b383c
313c0073
700f09db
623c1c73
38c3708c
55946007
0af209c3
301c0116
311c0b84
6c0c0000
36640cc6
500c8056
111c2046
21a30800
289b253c
32c3500f
011c0006
30830100
323c68d2
36e4164b
32c30494
700f7f72
32c3500c
011c0006
30830020
323c68d2
36e4158b
32c30494
700f7f92
32c3500c
011c0006
30838000
16546007
363c32c3
7872165b
100c700f
f88c103c
0080293c
280c313c
21e3a980
323c30c3
700f0fdb
27f21ac3
32c30f93
159b363c
fd737572
280c363c
0e73fd80
7492700c
277213c3
2a1b153c
313c300f
60070024
313c1e54
63d207c4
14946207
60073ac3
103c1654
700c0340
139b363c
74726d72
4bc3700f
6a548007
108c313c
784e69c3
2ac30cb3
363c44d2
fd80280c
400631c3
0001211c
69d23283
313c300c
