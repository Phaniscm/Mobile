681a4b2d
d51b07d2
07836818
492bd518
0158680b
2100d507
4106f2c2
46856808
be28f001
680ae00c
d4050251
f2c22100
68084106
e0034700
00e0f240
47086801
6801481e
d504028a
f2c22004
68014006
6803e00a
d50902db
5080f248
4004f2c2
f3c16801
02d13207
e004468d
6040f45f
4006f2c2
4a124685
01c06810
f04fd518
f1a3438c
f44f609a
60192100
f44f2201
234e0170
60416002
480a6043
01516802
6801d5fb
d5fc008a
f44f4b07
60182000
be3ef001
bf00e7fe
1208001c
24048580
24048604
46000058
46000004
00000000
00300920
003002e0
003003dc
0030040c
00300a94
0030098c
0030045c
003005e8
00300c0c
003008c8
00300488
00300684
00300274
003005a0
00300790
00300754
00300b3c
00300ba4
00300720
00300a88
003009ec
003006bc
00300c70
37300903
0000003d
0003e000
00437a31
40020000
00220000
007800d8
002000c7
00050001
00300fd5
00301075
00301099
003010c1
003010d9
003010f9
003011a9
00301265
003012a1
00301505
003015dd
00301691
00301105
00301715
003012dd
003056c9
00305cdd
00306889
00304669
00307947
00302051
00302061
003020c5
003020e9
00302105
00302135
00301f8d
00301fbb
0030215d
00301fa1
00301f8f
00302137
00301a6d
00301a83
00301d31
00301ac5
00304271
00304285
003036a5
00303b7f
00302259
00302417
003023d1
003023f7
00301919
003018e9
003011d9
003019f1
00300e91
00300ea3
00300f15
00300f39
00300fa7
00300fc7
00301a11
003015f9
00301aa5
00000004
0000000c
00000010
0000000c
00000014
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00302259
003024d3
003026a1
00303159
003031db
0030227d
003022c5
00303109
0030250d
003036a5
00303925
00302307
00303339
00303b7f
00302915
00302aa9
003038b1
00302441
00302469
003023d1
003023f7
00302417
00302881
00303ea1
00302385
00302ebd
00303315
00303f81
00303f91
00303f9d
00303fab
00303fb9
00303fd9
00303feb
00303ffd
0030400f
00304021
00304033
00304045
00304057
00304069
0030407b
0030408d
0030409b
003040ab
003040bb
003040cb
003040db
003040eb
003040fd
00304107
0030410f
0030411d
00304129
00304135
00304143
00304153
00304163
00304173
00304185
00304197
003041a9
003041bb
003041cd
003041df
003041f1
00304203
0030420f
00304221
00304233
0030423f
0030424f
0030425f
0030435d
00304271
00304285
00304299
003042ad
003042b9
003042d3
003042eb
00304305
0030431f
00304339
0030434d
003043b9
00304405
0030444d
0030449d
003044ed
0030453d
00304557
00304571
0030458b
003045a5
003045bf
003045d1
003045e9
00304615
00304641
00304669
00304657
003046b9
0030492d
003046c1
003046cd
003046d9
003046e1
00304963
003046f9
003046ff
00304985
003048dd
00304705
003049a5
00304895
00304919
00304923
00304d29
00304e5d
00304a53
003046bd
00304f27
0030525d
0030500d
00304f11
00304f2d
00305029
003052a7
00305487
003051fd
00305287
00305241
00306161
0030617d
003056c9
00305649
00305631
00306199
00305801
003061b5
00305811
00305821
003061d1
003061ed
00306209
00305831
00305849
003058c5
00305875
00305859
00305a3d
00306225
00306241
00305a4d
00305b09
00305a99
0030625d
00305a5d
00305a6d
00305a7d
00305c31
00305c3d
00305c49
00305c55
00305c61
00305c6d
00305c79
00305ccd
0030694d
00306b45
00305cdd
00306889
003062bb
00305d75
00306279
003067db
00305d9f
00306435
00306741
003066c5
00306651
003065dd
00305dc9
00306a09
003065bb
0030646f
00305df3
00305e05
00305e41
00305e53
00305e65
00305e77
00305e89
00305eab
00306561
00305f55
00305ef1
00306589
003064dd
00305fd5
0030603d
003060c7
00306bb9
00306bbd
00306bc9
00306bcd
00306bd1
00306bd5
00306bd9
00306be5
00306bf3
00306bf7
00306bfb
00306c01
00306c07
00306c0b
00306c0f
00306c13
00306bc1
00306bc5
00307311
00307219
00307189
00306d25
00306d35
00306ee5
00306f09
00306f15
00306ff9
00307165
00307175
00306c19
00306c25
00306c31
00306c3d
00306c49
00306c51
00306c5d
00306c63
00306c6f
00306c7b
00306c85
00306c91
00306c95
00306c99
00306c9f
00306cab
00306cb7
00306cc3
00306ccf
00306cdb
00306ce7
00306cf3
00306cff
00306d0b
00306d17
00301a6d
00301b1d
00301a51
00307325
00307c7f
00307351
00307361
00307bc7
00307add
00307a03
00307947
0030786d
00307d37
00307e13
00307373
003073a3
003076c9
00307ecd
00307eff
00307f03
00307f0b
00307f15
00307f19
00307f1d
00307f21
00307f2b
00307f35
00307f3b
00308561
00307f3f
00307f43
00307f47
003086e5
00307f4b
00308579
00308227
0030823d
00308523
003087b9
003083df
0030853d
003083e3
0030880d
00308813
00308817
0030881d
0030882d
0030883b
003088a1
00308853
003088e5
0030886f
0030888f
00308895
0030889d
0030890b
00308915
0030891f
0030892d
00308933
0030893b
00308945
0030894f
00308959
00308963
0030896d
00308a31
00308a81
00308979
003089d5
0030a21d
0030a25d
0030a2a1
0030a2e5
0030a329
0030a36d
0030a3e1
0030a469
0030a4ad
0030a535
0030a425
0030a579
0030a5b9
0030a059
0030a09d
0030a0e1
0030a125
0030a199
00309549
00308fa5
0030900d
003095ad
00309611
00308c51
00309679
003096e1
00309075
003090dd
0030994d
00308ab9
003099b1
00308cb9
00309a19
00309a81
00309145
003091ad
00309ae9
00309bb5
00308d21
00309b4d
00309c1d
00308d85
00309c85
00309ce9
00308de9
00309d51
0030a1dd
00308e4d
00309db5
00309215
00309265
00309e01
00309e4d
00309e99
00309f11
003094cd
00308e99
00309f89
00308ea1
00309ff1
00308ea9
003092b5
00308eb1
0030933d
00308eb9
00308ed1
003097b1
00308ee9
003093a9
00309745
00308f25
0030981d
0030988d
00308f05
003098b5
00309435
003098dd
0000ffff
0030a925
0030a5fd
0030a62f
0030a64b
0030a651
0030a663
0030a675
0030a67b
0030a693
0030a80b
0030aa3d
0030aabd
0030a817
0030a84b
0030a86d
0030a947
0030a8a5
0030abb1
0030ac55
0030ab15
0030a8c1
0030a8f9
0030ad63
0030ad67
0030afe1
0030afbb
0030af89
0030ae61
0030af0b
0030b029
0030b04f
0030b391
0030b075
0030aeef
0030b4d1
0030ad6b
0030ad71
0030ad81
0030ae29
0030ae1f
0030ad91
0030adaf
0030adb7
0030adbf
0030add3
0030adf1
0030ae0d
0030ae35
0030ae59
0030b7c5
0030b7c9
0030bed3
0030bea9
0030b885
0030b8a1
0030b7d7
0030b7e7
0030b7f7
0030b809
0030b81b
0030b82d
0030b83f
0030b84d
0030b859
0030b863
0030b7cd
0030b8bd
0030ba6d
0030bd61
0030bc1d
0030befd
0030c075
0030bc11
0030c4df
0030c493
0030c213
0030c25f
0030c2ab
0030c317
0030c33f
0030c367
0030c3a3
0030c52b
0030c52f
0030c533
0030c537
0030c53f
0030c547
0030c54d
0030c58d
0030c59d
0030c5ad
0030c5c5
0030c5dd
0030c5e3
0030c5e9
0030c5ff
0030c615
0030c61b
0030c621
0030c63d
0030c659
0030c661
0030c669
0030c66d
0030c671
0030c689
0030c69f
0030c6b3
0030c713
0030c73b
0030c745
0030c7d9
0030c7f7
0030c7fd
0030c9f5
0030c811
0030c815
0030c819
0030c821
0030c82f
0030c83d
0030c84b
0030c859
0030c86f
0030c885
0030c89b
0030c8b1
0030c8b9
0030c8c1
0030c8c9
0030c8d5
0030c8e1
0030c8ed
0030c8f9
0030c927
0030c92f
0030ca11
0030ca2f
0030ca4d
0030c94b
0030ca6f
0030c955
0030c969
0030c971
0030c979
0030ca91
0030cad3
0030c97f
0030c997
0030c9af
0030c9d3
0030c9c7
0030cb15
0030cbcf
0030cc0d
0030c9dd
0030ccb1
0030cf55
0030ccb5
0030ccbb
0030ccc1
0030ccd7
0030cced
0030ccf9
0030cd05
0030cd11
0030cd15
0030cd1b
0030cd1f
0030cd23
0030cd27
0030cd2b
0030ce11
0030cf71
0030cfb5
0030ce1d
0030ce4d
0030cf39
0030d059
0030d111
0030cfe5
0000ffff
0030d18d
0030d191
0030d197
0030d19d
0030d1b3
0030d1c9
0030d1df
0030d1f5
0030d20b
0030d20f
0030d213
0030d217
0030d21b
0030d21f
0030d419
0030d4a5
0030d2ff
0030d3fb
0030d561
0030d5e5
0030d4f9
03020100
00000000
01000900
00000302
09000000
0030d659
0030d65d
0030d663
0030d66b
0030d785
0030d673
0030d67d
0030da3b
0030d69f
0030d68d
0030d741
0030d73d
0030da75
0030da9f
0030dacb
0030d693
0030d777
0030d687
0030d699
0030d825
0030d8ed
0030da11
0030d745
0030d753
0030d765
0030db1d
0030dbf5
0030e30d
0030e235
0030e1a5
0030dc01
0030ddb7
0030df75
0030e757
0030e547
0030e747
0030e6bb
0030df91
0030e3e5
0030e42d
0030e4e5
0030ea1d
0030ea3d
0030ea59
0030e771
0030e7bf
0030e7f1
0030e829
0030eb71
0030eb89
0030ebc1
0030ebfd
0030ec2d
0030ec4d
0030ec6d
0030edc9
0030ea91
0030eac3
0030eae7
0030eb0b
0030eb3d
0030eb57
0030ef07
0030ef19
0030ef3b
0030ef4f
0030e931
0030e9f1
0030e9fd
0030e971
0030e979
0030e889
206e490a
20746567
20787220
2c746b70
42207852
65666675
6e692072
20787220
20616d64
63736564
20736920
4c4c554e
490a000a
7573206e
74696d62
20787220
20746b70
5852202c
66756220
20726566
61207369
6165726c
76207964
64696c61
490a000a
7573206e
74696d62
20787220
20746b70
5852202c
66756220
20726566
6e207369
6120746f
6c696176
656c6261
200a000a
65636572
5f657669
6d6f7266
5f61745f
656e6f64
7273695f
6552202c
76696563
4e206465
204c4c55
6b636150
0a207465
344d0a00
52534920
75202c20
7078656e
65746365
6e692064
72726574
20747075
0a000a20
66206e49
656d6172
69727720
2c206574
766e4920
64696c61
20585420
6d617266
65642065
69726373
726f7470
0000000a
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
2300b510
d0034293
54c45ccc
e7f93301
b510bd10
18424603
2c3f1ad4
2400d912
605c601c
60dc609c
615c611c
61dc619c
625c621c
62dc629c
635c631c
63dc639c
e7e83340
033ff021
f00118c0
4603043f
1ad21902
d9062a0f
601a2200
609a605a
331060da
f004e7f4
19000430
010ff001
18424603
2a031ad2
2200d903
2b04f843
bd10e7f7
f021b570
f0010503
46290403
f7ff4606
b134ffbe
19041970
f8002300
42a03b01
bd70d1fa
0303f022
47f0e92d
0c03eb01
425b18c6
0503eb0c
351018f4
f1133410
da110f0f
ac0cf855
9c08f855
8c04f855
7c10f855
ac0cf844
7c10f844
9c08f844
8c04f844
e7e83310
0f03f113
f85cda04
50f44003
e7f73304
0303f012
1ad2d007
18891880
e8bd461a
f7ff47f0
e8bdbf77
b53087f0
5cc52300
42a55ccc
d806d305
429a3301
2000d1f7
2002bd30
2001bd30
b122bd30
f8001882
42901b01
4770d1fb
f8d04b23
681a14c8
34c4f8d0
41f0e92d
f8d24604
f50050cc
18c970ea
723af44f
f89447a8
b9100496
f8842201
7a632496
1496f894
0020f003
b33ab2c2
252c4f14
76eaf504
6839434d
0805eb06
64a9f504
46206b0b
59724798
f8d86838
f8d03004
18d3c0a4
5090f04f
47e02100
4809683a
30ccf8d2
220c4621
59714798
60014806
2004f8d8
48055973
600118d1
81f0e8bd
24060ff0
24060030
24060028
2406002c
88134a06
512cf423
0c59044b
4020f440
80114b03
801ab282
bf004770
4105003c
41050034
88134a08
402bf403
d0f92800
88138811
502cf423
0c580443
f4218010
0451522c
47700c48
4105003c
60184b04
22013308
6818601a
d5fc0702
bf004770
4600816c
68194b04
d0034208
4b044a03
60186010
bf004770
4105008c
46008180
41050090
60184b01
bf004770
41050090
4b24b538
f012681a
46057280
f04fd011
22015190
212cf8c1
5390f04f
012cf8d3
d4f907c0
20c4f8d3
1104f042
10c4f8c3
4819e026
68014c19
0f01f011
6803d00a
d5070799
49166820
30a8f8d0
5090f04f
e0154798
20016822
478868d1
68436820
47982056
68114a0d
47806888
d10528bb
681a4b08
7180f042
e0016019
d1f128dd
68184b06
f8d04629
f04f20ac
47905090
bf00bd38
24048580
1208001c
24060ff0
2406003c
f890b508
b9133496
f8802301
212c3496
0303fb01
f8d34a05
f8d011d4
681204c4
f8d21840
304020b8
bd084790
24060ff0
4b20b5f0
68184606
2240b093
40ccf8d0
a8024631
f8bd47a0
f6452008
428a21a5
f8bdd12e
2300500a
ac124f16
1c5f6838
01c3eb04
04c7eb04
30ccf8d0
2c40f854
0c34f851
427ff022
479819a9
0c40f854
2c3df814
0117f3c0
440d09d2
d0e3463b
49099803
20b8f8d0
92006008
30c0f8d0
99019301
f8d04668
4708d000
bdf0b013
bf00e7fe
24060ff0
e000ed08
4d0db570
f5004606
cd0f74dc
e895c40f
e8840007
7a330007
0040f003
b149b2c1
f8968932
f3c211be
1c5813c1
0102f360
11bef886
bf00bd70
00300134
4607b5f0
460eb087
490bb1a2
f8d06808
92015098
24009a0c
bf082b02
93002303
71dcf502
94039402
f04f9404
463a5090
47a84633
bdf0b007
24060ff0
b5706a0b
0399460c
46154606
6a10d410
d50d0382
680a4983
005cf104
30ccf8d2
015cf105
47982204
f4406a20
62213100
03536a22
6a2bd410
d50d0358
68014879
f8d12206
f10430cc
f1050060
47980160
f4426a22
62202080
03096a21
6a2bd410
d50d031a
68104a6f
0166f105
30ccf8d0
f1042204
47980066
f4416a21
62222200
06036a28
68a9d517
68ea686b
60a16928
606369a9
696b60e2
612069ea
6a2061a1
1554f8d6
61e26163
0380f040
0280f021
f8c66223
f8d42554
07583090
f8d5d407
07410090
f043bf44
f8c40304
f8d43090
050a1094
f8d5d409
05102094
6fabd505
6000f441
f8c467a3
f8d40094
05593094
f8d5d409
054a1094
6fead505
6080f443
f8c467e2
f8d40094
06983090
f8d5d40b
06891090
f8d5d507
f04320ac
f8c40020
f8c420ac
f8d40090
065a3090
f8d5d40b
06481090
f8d5d507
f04320b0
f8c40040
f8c420b0
f8d40090
04d93090
f8d5d413
04ca1090
4a33d50f
f1056810
f8d001e0
220c30cc
00e0f104
f8d44798
f4411090
f8c45280
f8d42090
06030094
f8d5d413
06183094
4927d50f
f504680a
f8d27096
f50530cc
221c7196
f8d44798
f0400094
f8c40180
f8d41094
00d93090
f8d5d40b
00d22090
f8d5d507
f0430168
f8c45180
f8c40168
6a2b1090
d50b019b
6a206d6a
3554f8d6
f0406562
f0237100
62217200
2554f8c6
01406a28
6da9d50b
f8d66a23
65a10554
6280f043
6180f020
f8c66222
f8d41554
06993094
f8d5d40b
06922094
f8d5d507
f0431170
f8c40020
f8c40094
bd701170
24060ff0
47f3e92d
682b4d32
46049000
0628f100
f8d06a1f
22020530
46312301
f8b447b8
f6459028
4581205a
6829d14e
6a0f9400
0530f8d4
2300226c
47b84631
f104682a
6b57080c
46202301
46324641
682b47b8
20709400
f1046a1f
23020198
7290f44f
f8d447b8
048300b8
6829d524
a0b4f8d4
f5049400
220267ab
c020f8d1
46502301
47e04639
454a8d22
4b12d114
02006818
6829d510
f8d19400
f10ac020
1cb90002
72c7f44f
47e02301
4620682d
46316bab
4798463a
68104a06
6b454641
46204632
47a82300
e0002001
e8bd2000
bf0087fc
24060ff0
24048580
4c05b538
68196823
47884605
69826820
47904628
bf00bd38
24060ff0
7a06b5f7
31bff890
0683f3c6
1307f366
f8804605
460c31bf
6a40b141
491bb930
4630680a
70b4f8d2
47b82101
30b8f8d4
00c0f8d4
93004916
600c9001
f0027aea
b2fb0702
21ecb143
46202201
f9e4f000
70ecf8d4
e00342b8
70ecf8d4
4287480d
2700bf14
b13c2701
b9296a69
68134a07
f8d34630
479020b4
9901b12f
f8d4466c
4708d000
2001e7fe
bf00bdfe
24060ff0
e000ed08
10ad10ad
4d1fb5f7
4604682b
478869d9
f8947a26
f3c601bf
f3660683
f8841007
682a01bf
f8d22000
47b870bc
4630682b
20b4f8d3
47902101
46306829
70b0f8d1
47b82100
27006828
f8d09700
2201c09c
5090f04f
f504463b
47e071dc
f8c4682b
6a5a7530
47904620
2001b110
62606120
46046829
30b4f8d1
21004630
46204798
bf00bdfe
24060ff0
461fb5f7
46146a13
4606039a
d523460d
0554f8d0
3300f410
4a68d11e
1080f8d2
1186f363
1080f8c2
0080f8d2
0380f040
3080f8c2
408cf04f
06936d82
4960d5fa
f8d14b60
f8b4e000
f8b4205e
f8de105c
4359c03c
47e0435a
01406a20
f8d6d50d
f0122554
d1086280
48574955
2101680b
c04cf8d3
3074f895
6a2047e0
d5120181
2554f8d6
7100f012
4b4dd10d
681a484d
fbb36f2b
2001f3f0
f8d29000
484bc048
460bb29a
6a2147e0
d50d034a
2554f8d6
d4090353
f8944b42
68181060
2062f8b4
f04f6c03
4798408c
03086a21
f8d6d514
03112554
483ad410
e069f894
f8cd6800
f8d0e000
f894c044
f8941066
f8942067
f04f3068
47e0408c
061a6a23
f8d6d52a
060b1554
7a62d426
0080f002
b143b2c3
f89568a1
f3c101b2
f3624202
f8850002
686301b2
31acf8c5
f50568e2
608a71d6
60c86920
610b6963
4b2169a2
69e0614a
6188681a
93002300
c09cf8d2
5090f04f
47e02201
b1176a21
1554f8c6
0608e02d
6868d51a
f040491a
606b0302
2088f894
0080f8d4
616860aa
0a9a680b
d50a0751
0303f002
fa012120
b2d3f203
bf944298
60eb60e8
60e8e000
0090f8d4
d50c00c2
f8d54907
680b24b8
1168f8d4
30ccf8d3
f2051889
226040c4
bdfe4798
24048400
24060ff0
000f4240
24041400
24042000
2404860c
bf9a2804
5c1b4b09
f1032300
f503538c
00835080
f022681a
601800c0
6819b121
0280f041
4770601a
bf004770
0030012c
41f0e92d
280d4606
e8dfd829
2c07f000
28100a0d
2c072828
1310280d
24002501
2502e023
e0202434
242e250a
2502e01d
e01a243a
49244b23
601a2201
20004b23
60082208
60886048
610860c8
61886148
620861c8
62886248
e8bd601a
240081f0
46262501
250ae001
b1192406
d8162e04
81f0e8bd
eb07460f
fa5f0804
2100f888
46424813
f002462b
4812fb84
37016801
2094f8d1
47904640
d1ec2f06
2434e7e6
46222100
480a230a
fb73f002
68184b09
1094f8d0
34014620
4788b2e4
d1ef2c3a
81f0e8bd
460081b4
46006000
460081c0
46130000
24060ff0
2801b138
f04fd10b
f44f438c
601a2280
f04fe005
f44f418c
608850c0
47704770
b1d1b530
0503f021
42ab2300
58c4d205
bf281912
33043201
f011e7f7
d00a0103
f04f00c9
58c334ff
f101fa04
0001ea23
bf281882
43d03201
4610bd30
0000bd30
681a4b05
d5010711
bb1ef7ff
60182001
070a6819
e7f7d5fc
46008174
f7ffb508
f7fffb01
2831fb11
38aad0fb
2001bf18
b940bd08
00b8f240
468d6801
00c0f240
47086801
28014770
f240d103
680100e0
47704708
210cb508
6300f04f
34c4f8c0
f500460a
f7ff60a9
e8bdfa86
f0024008
0000b965
681a4b08
0001f042
60184a07
f4416811
60101000
07d0681a
6819d5fc
dafc2900
bf004770
20280014
46008044
698bb508
f8d1b17b
f01330b0
d00a0380
0180eb01
3148f8d1
4610b12b
30004798
2001bf18
4618bd08
0000bd08
4c4eb538
68252b01
4b4dd167
60186824
6000f04f
88016219
f645625a
4291225a
f8d0d115
049a3090
f8d0d509
180a108c
6a10d005
d5020603
1d114842
f04fe009
6a196300
d5020608
493f483e
483de001
221c493e
f9e2f7ff
48394a3c
60836853
11c1f3c4
1c4b7a82
0202f363
72827ac3
0140f3c4
0283f3c4
03c3f361
1307f362
2407f3c4
f00472c3
b2dc0320
f04fb304
f8d25290
f8d21100
628130fc
f8d262c3
f8d210d8
630130dc
f8d26343
4b2810e0
68196381
d40b01c9
30c8f8d2
10ccf8d2
f8d263c3
f8d230d0
640120d4
64826443
68184b1f
6080f040
2b02e02d
4b1cd10f
f442681a
601a1200
b1084b15
e0016058
60584818
bf082900
60994619
2b03bd38
4b0fd102
bd386019
d1042b04
68194b10
0080f441
2b05e00f
4b0dd10e
f422681a
6019217f
f3c0681a
ea4220c7
60193100
f442681a
60181080
bf00bd38
24048604
24060000
24060004
08000004
00300134
24048580
24060c00
4b25b5f7
48264c25
f8d0681e
602010bc
47882000
f3c66822
f8d20583
462870b4
47b82101
46286823
20b0f8d3
47902100
68202500
22019500
709cf8d0
f04f4919
462b5090
682147b8
2607f3c6
308cf8d1
f0064798
b2d60220
6820b176
48126b01
4b124788
681a6824
40a4f8d4
46291d18
f04f6803
47a05090
480e490d
f022680a
600b6380
68014a0c
20206011
4006f2c2
47086801
bf00bdfe
24048604
24060ff0
00300150
24060004
24060030
24060028
24048580
24060024
e000ed08
681a4b8b
b57002d0
681ed509
f3c66819
02d03207
5480f5a0
1580f421
6818e008
f4104c84
d0041f00
68a46819
1500f421
4620601d
61ddf44f
f8d4f7ff
4b7c4e7e
681d487e
68016832
60254e7d
606260a1
4b7c6832
07d14d7c
d404602b
6801487b
d40007ca
f8d3e7fe
462030e0
7a254798
0602f005
2a00b2f2
8090f000
68304e72
108cf8d0
68334788
6add4620
280047a8
6a60d07c
050cf104
d04a2800
1500f8d4
33bbf64b
d1184299
20004629
f7ff4622
4601fe87
f0402800
683080b2
2504f8d4
32406f03
47984620
46292001
f7ff4622
2800fe77
80a3f040
2002e00d
46224629
fe6ef7ff
f0402800
f8d4809a
f02220b8
f8c40620
f8d460b8
485320b8
0f20f012
f8d4bf1c
600110d4
d50804d6
220c6801
60ccf8d1
60a9f504
7184f504
f8d447b0
065830b8
f8d4bf4c
f44f30d8
f8c43380
f8d434c8
075120b8
4845d504
f0416801
60060601
4e407ae3
0250f003
d10b2a40
46292003
f7ff4622
2800fe33
6830d15f
46206a86
e7fe47b0
46292004
f7ff4622
2800fe27
6835d153
1198f8d4
34c4f8d4
20dcf8d5
18c94620
e0484790
f8d46832
f8d214c4
462060dc
e04047b0
f0007ae0
b2cb0140
4e26b303
68324d27
0001f012
f8c4d106
682c0538
2084f8d4
e7fe4790
68c16828
47882001
689e682b
682a47b0
f8d22033
47881080
682dbb08
0538f8c4
6084f8d5
e01a47b0
0504f000
b1b6b2ee
0208f000
b930b2d0
4e164913
f8d3680b
47a8508c
4e14e000
f64a6832
428220bb
490dd105
680b68b0
50b8f8d3
4d0a47a8
46206829
30dcf8d1
47982100
bf00e7fe
24048580
24060000
24048584
24048604
1208001c
00300150
24060ff0
46008010
24048600
0017fff0
0030fff0
b11ae7fe
d1032a01
47708001
47707001
47706001
b119b082
d1032901
e0028803
e0007803
93016803
b0029801
e92d4770
9e0743f0
d90642b3
d1062b02
bf0c2e00
27022704
2701e002
2702e000
2400b3c2
462546bc
d00f2e01
2e02d304
6805d115
e0122404
9000f814
08c4ea4f
f808fa09
0508ea45
e0083401
9000f834
08c4ea4f
f808fa09
0508ea45
f1bc3402
d1e10c01
19001b12
d0d92c00
d0082b01
2b02d302
e00cd00a
5b01f801
0a2d3c01
f821e7f2
3c025b02
e7ed0c2d
5b04f841
e7fee7c6
83f0e8bd
08988803
f110bf00
d2fb30ff
00004770
b5f74603
6899460c
6840681b
b29a4d14
32010e1e
0f01f016
f026d118
f006067f
b12e07ff
61bdf894
0601f046
61bdf884
9400682d
f3c36a2d
47a85381
f894b177
f36f01bd
f8840000
e00701bd
f3c3682c
95005501
f3c36ee4
47a05381
bf00bdfe
24060ff0
4604b510
78a14b06
f3c16818
6f421101
47906860
68e168a3
42884018
bd10d1f2
24060ff0
4a05b510
68114603
6f8c7882
68996840
47a00992
bf00bd10
24060ff0
4d0ab538
682b7881
6f5a4604
f3c16880
47901101
78a26861
68284001
6f836925
432968e0
47980992
bf00bd38
24060ff0
b0824770
78cb9201
d40b07da
0102f003
b102b2ca
f8c02201
f8d02534
b1080534
47089901
4770b002
4605b5f0
b111b089
93028d43
9202e000
68014838
6a0c9500
22049802
a9032302
f89d47a0
4b34200e
053cf8d5
060ff002
6026f853
f89db130
f001100f
b2d30220
d0352b00
000ff89d
0140f000
2a00b2ca
4c28d02e
68279b02
1d189500
6a3fa904
23021f32
f89d47b8
f000000e
2905010f
e8dfd81b
0603f001
1714110c
6d036820
6823e007
6d5aa803
47904629
6822e010
a8036d93
e00b4798
6dcb6821
6820e7f9
e7f66e03
6e536822
6821e7f3
47986e8b
100ff89d
0206f001
d10a2a02
f8d5480d
680320a4
01a0f105
46286fdb
b0094798
9c02bdf0
f0011930
b2f30608
2b009002
4904d096
9500680a
a9026a14
23022204
e78d47a0
24060ff0
00300234
1080f8c0
69016402
400a4a05
0102f042
3343ea41
6a026103
d4fc07d3
bf004770
ffdf9ff8
4604b5f8
460f4615
2108461e
463a462b
ffe4f7ff
7a706923
f000490a
40190280
010cf041
2b00b2d3
f44fbf14
20001000
3545ea41
61254305
06126a22
6c23d4fc
bdf8b2d8
07c78000
4604b5f8
4616460f
22062108
f7ff461d
6920ffc1
51fff420
021ff021
0301f042
46206123
ea462110
462b2207
ffb2f7ff
f4206920
f02151ff
f042021f
61230301
b570bdf8
9d059c04
f101b910
e0016100
6110f101
fbb41c58
fb00f6f0
b10e4616
1ba41824
1914b94b
42a34613
1a98d004
f8035c40
e7f80b01
2b01bd70
4613d10e
42831910
8808d009
0b02f823
07c07ba8
3101d501
3102e7f4
bd70e7f2
d10d2b03
19104613
d0094283
f8436808
7ba80b04
d50107c0
e7f43102
e7f23104
0000bd70
681a4b0f
0220f042
7900601a
1240f3c0
f0400210
f442528d
60082046
bf00220a
d1fc3a01
f0206818
601a0220
4b056808
600b4003
4804680a
0300ea42
4770600b
460081bc
01ac6100
01ac6101
f8c0680b
684a30c8
20ccf8c0
f8c0688b
68c930d0
10d4f8c0
20c4f8d0
0304f042
30c4f8c0
680b4770
30d8f8c0
f8c0684a
688920dc
10e0f8c0
30c4f8d0
0202f043
20c4f8c0
b5304770
50c4f8d0
5480f44f
f401fa04
f8c0432c
f1c140c4
f1c1043f
eb00013e
eb000484
60620081
bd306043
21004602
4807b508
f8b9f002
21004805
f874f002
21004803
f8baf002
d0f92800
bf00bd08
24042000
43f8e92d
46154604
22064689
46982108
9f08462b
feecf7ff
f4266926
f02050ff
f041011f
61220201
21084620
462b2242
fedef7ff
45462600
4620d007
464a2108
f7ff462b
3601fed5
6923e7f5
50fff423
011ff020
0201f041
b1276122
e8bd4638
f7ff43f8
e8bdbfb9
690383f8
53fff423
031ef023
6103b510
6843b932
0206f023
0141ea42
bd106041
00533203
22036944
f203fa02
0202ea24
f103fa01
61414311
0000bd10
43f7e92d
790e6903
f423460c
461751ff
021ff021
0301f042
78216103
0641f3c6
f0014632
46050103
ffcdf7ff
f8947a20
78a38000
0202f000
f008b2d2
b13a0803
f3c28922
46280287
ea422110
e00a2203
f00179a1
28010007
f407bf04
00d27280
21084628
4633431a
fe70f7ff
f3c37823
45410181
4628d007
f7ff4632
f894ffa4
f3ccc000
79a10881
d003074a
0007f001
e00000c1
463a2108
46284633
fe56f7ff
f0027862
b2d90310
f002b189
45410103
4628d007
f7ff4632
f894ff86
f0088001
46280803
22002108
f7ff4633
78e0fe3f
0ff0f010
89e2d104
63f0f402
d04c2b00
78e189e7
f3c77823
010210c3
1711ea42
45410999
4628d007
f7ff4632
f894ff64
ea4fc000
7861189c
0008f001
bb2ab2c2
05b87a63
027ff023
01fff002
69280d83
4a1bb122
f4424002
e0011220
40024a18
0004f042
3246ea40
03c3ea42
ea430ab8
612a62c0
061b6a2b
6c28d4fc
b282b109
b2c2e000
92013f01
e00ed1f4
0903f017
f04fbf08
46280904
ea4f2200
463301c9
fdecf7ff
0709ebb7
7821d1f0
1101f3c1
d0034541
46324628
ff1df7ff
83fee8bd
07c78000
4ff7e92d
78cf790e
0641f3c6
46044692
f007460d
8b4a070f
6843b91e
0841f3c3
6943e008
0803f106
0048ea4f
f100fa23
0803f001
10c4f8d4
f0117ca8
f0000f08
f04f0307
d00e0901
d8042b03
fc03fa09
190cea4c
1f18e009
f300fa09
1103ea43
2901ea4f
fa09e001
6920f903
53fff420
011ff023
0001f041
7a2b6120
0102f003
b128b2c8
0f03f1b8
2110d101
0a12e001
46202108
f7ff4633
2f09fd8f
f1b8d108
d1050f03
21204620
46332200
fd84f7ff
0202f1a8
d90e2a01
07db7bab
f8d4d520
f42110c4
f8c42000
210300c4
46324620
feaff7ff
8a6fe014
17c3f3c7
d0eb2f00
0b03f017
f04fbf08
46200b04
ea4f2200
463301cb
fd60f7ff
070bebb7
e7dbd1f0
0371792a
0206f002
f8d4b122
f4100094
e0033f00
3090f8d4
3f80f413
f8d4d103
071830c4
6920d50e
40034b2c
f0007a68
b2c00080
bf142800
1020f44f
f0432000
e00d0314
4b256920
7a684003
0080f000
2800b2c0
f44fbf14
20001000
030cf043
4303430b
6a236123
d4fc061b
f8d4b122
f4133094
e0033f00
0090f8d4
3f80f410
f8d4d103
070000c4
6c23d502
e001b298
b2d86c23
98019001
0f00ea19
7baad1b4
d50507d1
10c4f8d4
2300f441
30c4f8c4
46414620
f7ff4632
6920fe3c
52fff420
011ff022
0301f041
f1ba6123
d0020f00
f7ff4650
9801fde5
8ffee8bd
07c78000
43f8e92d
f8bd9d09
46068020
4691460c
b90d461f
e000684b
2108694b
46202206
f7ff462b
6921fcd9
50fff421
021ff020
0301f042
61232108
464a4620
f7ff462b
78f1fccb
020ff001
46202a09
2120d101
2108e000
462b463a
fcbef7ff
46202108
462b4642
fcb8f7ff
f4206920
f02353ff
f041011f
61220201
f00078f0
2b0a030f
4620d106
22004631
43f8e8bd
bec8f7ff
83f8e8bd
4ff8e92d
6843469a
f891790e
f8ddb003
f0139028
46040840
4617460d
0641f3c6
0b0ff00b
6840d008
0140f020
6a226061
d4fc04d0
0801f04f
f0037beb
b2c10010
f8d4b129
f4222130
f8c45380
7ba83130
d50507c1
10c4f8d4
2200f441
20c4f8c4
46207aeb
0103f003
f7ff4632
f1b9fda8
d1050f00
f0037a6b
b2c10080
e012b941
f0206920
61217100
04526a22
e7f1d4fc
0f09f1bb
d1034620
f2402110
e01062f9
22062108
4620e00d
46332206
f7ff2108
7a2afc49
0302f002
b128b2d8
21084620
463322f9
fc3ef7ff
f4216921
f02353ff
f040001f
61210101
f0037a2b
b2c10002
bf0c2900
21102108
d1012f20
e0038aea
bf0c2fd8
8aaa8a2a
46334620
fc22f7ff
d00c2fc7
075379aa
f002d003
00d90307
2108e000
46524620
f7ff4633
6920fc13
51fff420
021ff021
0301f042
46206123
9a0b4629
fe2af7ff
07c07ba8
f8d4d505
f42110c4
f8c42200
f1b920c4
d1030f00
0f01f1b8
e007d10f
f0436923
61207000
04496a21
e7f3d5fc
f0426862
60630340
04c26a20
7be9d5fc
0210f001
b90bb2d3
8ff8e8bd
0130f8d4
5180f440
1130f8c4
8ff8e8bd
4ff0e92d
b08b460d
f8bd79aa
792e1058
46989102
f8dd78eb
f0029050
46040107
f0032904
f3c6000f
90010641
00c8d006
fa022201
1e4bf100
0803ea08
f0106860
d0090240
f0216861
60630340
04c26a20
2201d4fc
e0009207
7be99207
0310f001
b128b2d8
2130f8d4
5180f422
1130f8c4
07db7bab
f8d4d505
f44000c4
f8c42200
210020c4
f8dd2301
f8cda054
f8cd9014
f8cd9010
46c3900c
93069100
0f00f1ba
8138f000
46207aef
0103f007
f7ff4632
7a68fcbc
0280f000
b151b2d1
2a099a01
d1034620
f5022110
e01062de
22062108
4620e00d
21084633
f7ff2206
7a2bfb69
0702f003
b128b2f8
21084620
463322f9
fb5ef7ff
f4216921
f02353ff
f047071f
61200001
f0027a6a
b2cb0180
b15b7aaa
29099901
7b2bd105
21104620
2202ea43
4620e00f
e00c2108
21084620
f7ff4633
7a2ffb3f
0002f007
b12ab2c2
46207b2a
46332108
fb34f7ff
b1cf9f06
46207aea
0181f3c2
f7ff4632
79a9fc68
d0030748
0007f001
e00000c1
46332108
465a4620
fb1ef7ff
f1b37aab
bf1807af
97062701
07d27baa
f8d4d50c
f42110c4
f8c42000
7aeb00c4
1201f3c3
0730f043
72ef9200
1e489902
0300ea1b
9a02bf1b
0302ebc3
b29b460b
bf284553
b29f4653
0a0aebc7
2f0044bb
7ae9d067
f3c14620
46321101
fc2bf7ff
6960796b
0140f3c3
020ff020
f106fa01
61614311
f0007be8
b2d90320
9917b339
981b4a86
1080f8c4
b1a86122
2115981c
fd18f001
f001981c
981cfd05
f0012115
2800fe52
f5a7d0f9
46207780
46324629
f7ffb2bf
e7cafce7
991b981d
fad5f002
2100981d
faaef002
d1f92800
9a17e7eb
9b03b952
2b01f813
93034620
46332108
faacf7ff
e01a3f01
28019817
9b04d10a
2b02f833
93044620
46332110
fa9ef7ff
e00c3f02
2b039b17
9b05d1a1
2b04f853
93054620
46332120
fa90f7ff
b2bf3f04
9a18e795
7baab99a
d51807d3
10c4f8d4
f4419a00
f8c42000
7aeb00c4
1305f362
72eb4611
46324620
fbb5f7ff
6921e007
7000f021
6a236120
d4fc0458
6961e7e3
000ff021
782b6160
f0034620
46320103
fba1f7ff
46204632
f7ff4629
9a19fc83
4610b112
fb4ef7ff
29009918
aeccf43f
f0406920
61237300
04516a22
e6c3d5fc
f0007a68
b2d10280
9901b151
46202909
2110d103
42fbf240
2108e010
e00d2204
22044620
21084633
fa38f7ff
f0037a2b
b2c20002
4620b12a
22fb2108
f7ff4633
6923fa2d
50fff423
021ff020
0101f042
7bab6121
d50507da
00c4f8d4
2200f420
20c4f8c4
29019907
7be9d00b
0310f001
b170b2d8
2130f8d4
5180f442
1130f8c4
6863e007
0040f043
6a226060
d5fc04d3
9b1ae7eb
f1b4b35b
d1025f80
6080f04f
f1b4e004
d1025f90
6000f04f
23009009
1ad29a15
d9092a03
eb089909
f8590001
58c01003
d1034288
e7f13304
e0012000
30fff04f
429318d2
9c09d00d
0104eb08
4003f819
428c5cc9
3301d103
981ae7f3
f04fe001
b00b30ff
8ff0e8bd
00200802
5f90f1b0
43f8e92d
4b8dbf0c
681e4b8d
070ff016
460d4604
1841f3c6
0980f006
4639d125
f7ff462a
4620faf6
22ff2108
f7ff462b
6923f9b3
50fff423
011ff020
0201f041
46206122
462a2102
fae3f7ff
21084620
462b22ff
f9a0f7ff
f4236923
f02050ff
f041011f
61220201
f1b9e0e0
d0070f00
f4436943
61603080
f4416961
61624200
46414620
f7ff462a
2f01fac4
80c3f000
d1122f02
21084620
462b22ff
f97cf7ff
f4236923
f02050ff
f041011f
61220201
21104620
72fff64f
2f03e004
4620d10e
22ff2108
f7ff462b
6923f967
50fff423
011ff020
0201f041
e09c6122
d1192f04
0f00f1b8
8097f000
21084620
462b22f5
f952f7ff
f4236923
f02050ff
f041011f
06f30201
d5016122
e0002096
f7ff2032
e080fa37
d10e2f05
21084620
462b2206
f93af7ff
f4236923
f02050ff
f041011f
61220201
2f06e7c3
f1b8d114
d06a0f00
21084620
462b2266
f926f7ff
f4236923
f02050ff
f041011f
61220201
21084620
e7c42299
d1162f07
0f00f1b8
4620d053
f2462110
462b6299
f90ef7ff
f4236923
f02050ff
f041011f
61220201
21104620
1266f649
2f08e7ab
2100d11c
460b220d
f0014828
2100f822
460b220d
f0004825
2100ff8f
220d4823
f000460b
06f0ff81
2096d501
2032e000
f9daf7ff
2100481d
e01d220d
d11e2f09
220e2100
4819460b
f803f001
220e2100
4816460b
ff70f000
220e2100
4813460b
ff62f000
d50106f1
e0002096
f7ff2032
480ef9bb
220e2100
f0002301
f1b9ff5d
d0070f00
f4236963
61603080
f4216961
61624200
21004620
e8bd462a
f7ff43f8
bf00b9ec
24048584
41300584
46130000
4615b570
2a059a04
460e4604
2a09d004
2238bf14
e0002200
2e022235
d1124620
462b2108
f894f7ff
f4236923
f02050ff
f041011f
61220201
46314620
e8bd462a
f7ff4070
4629b9c2
4070e8bd
beb2f7ff
41f0e92d
460e4604
461d4690
6842b91b
0741f3c2
6943e006
00781cef
f100fa23
0703f001
21084620
2206462b
f868f7ff
3008f898
0002f003
b139b2c1
d1052f03
21084620
462b22f9
f85af7ff
f4226922
f02353ff
f040001f
61210101
2e08b10e
4620d10d
22502108
f7ff462b
6922f849
53fff422
001ff023
0101f040
e8bd6121
e92d81f0
79164ff7
f3c678d7
46040641
4615468b
f0074698
b91e070f
f3c26842
e0080941
f1066943
ea4f0903
fa230049
f001f100
f1b80903
f8b50f00
da03a018
4800f028
e0002301
7ba82300
07c19301
f8d4d505
f44110c4
f8c42200
462020c4
462a4639
f7ff4633
2f08ff8b
2f03d001
4620d10d
22062108
f7ff4633
6923f801
50fff423
011ff020
0201f041
7a2b6122
0002f003
b131b2c1
0f03f1b9
2110d101
ea4fe002
21082a1a
46524620
f7fe4633
2f09ffe7
f1b9d109
d10c0f03
21204620
46332200
ffdcf7fe
2f03e005
2110d101
2f08e005
9a01d0fb
d1f82a00
792b2108
0f06f013
f8d4bf15
f8d43094
f3c33090
f3c34340
46204300
2110b11b
220bea4f
465ae000
f7fe4633
6920ffbb
51fff420
021ff021
0301f042
46426123
46294620
f9d2f7ff
07c27ba8
f8d4d505
f42110c4
f8c42200
e8bd20c4
00008ffe
5f90f1b0
4b05bf0c
681a4b05
003ff022
681a6018
60194311
bf004770
24048584
41300584
43f7e92d
4617780b
0230f003
f1b24605
f1d00020
f0030900
eb590803
f1b80900
460c0f03
f1b8d007
bf0c0f02
0804f04f
0800f04f
f04fe001
78e60808
060ff006
f2002e0a
e8df815d
000bf016
000b015b
001200e3
015b001b
00e300a6
0118004e
79227823
46289600
1101f3c3
f1b9e035
f0000f00
79238145
213e4628
e13b2280
96007923
f3c32100
46280241
f7ff460b
f1b9fe9f
d0160f00
463a4621
f7ff4628
7be2f963
0140f040
0040f002
b123b2c3
f0410209
f0470108
46284700
4622b289
f7ff463b
7822feee
0303f002
f0402b02
79228117
46289600
f3c24619
23000241
fe76f7ff
2a30e10c
f894d10d
f00cc009
fa5f0e80
f1b8f88e
bf0c0f00
0801f04f
0802f04f
f04fe001
79220800
21009600
4628460b
0241f3c2
fe5af7ff
78e189e6
10c3f3c6
ea43090b
2a081200
2a10d904
2602bf94
e0002600
7be02606
0140f000
b17bb2cb
463a4621
f7ff4628
0202f90d
417ff402
f0414628
4622010f
4300f047
fe9ff7ff
96007920
0341f3c0
46209301
22724629
7340f44f
f9e6f7ff
f8cd7922
f3c28000
91010141
46294620
23002272
f9daf7ff
7923e0b4
21009600
0241f3c3
460b4628
fe14f7ff
78237a66
f00678e1
b2c20004
00c0f003
bf0c2a00
22002208
ea4f2840
d1011611
e00400b6
d1012880
e0000076
796100f6
1302f3c1
7923431a
21814628
1206ea42
0341f3c3
fecef7fe
0f00f1b9
7822d107
0030f002
bf142810
229f22df
225fe000
46287923
e0732161
96007923
f3c32100
46280241
f7ff460b
4621fdd7
4628463a
f89ef7ff
0949ea4f
2000ea49
463bb281
46224628
fe31f7ff
f0017821
2b020303
7922d15a
46289600
f3c24619
23000241
fdbaf7ff
282f78e0
f000d906
293001f0
2230bf14
e0002220
46282200
230021c0
7a61e040
077ff021
f987fa5f
0f00f1b8
78e2d00e
03c0f003
ea4f2bc0
bf181012
28080040
2810d906
4607bf8c
e0022704
e0004647
79232700
21009600
0241f3c3
460b4628
fd88f7ff
79237961
1202f3c1
1042ea47
0141f3c3
9101b287
46209700
22714629
f7ff2303
f1b8f933
d1020f00
0f00f1b9
7923d008
21314628
0209ea48
0341f3c3
fe46f7fe
78227a61
0380f001
0003f002
2a00b2da
2104bf14
43012100
08c37ce0
1141ea43
b0034628
43f0e8bd
be58f7ff
a904b538
b189c932
46202114
f836f001
f0014620
4620f823
f0012114
4620f981
f0012114
2800f96c
bd38d0f9
f0014628
4628fdf8
f0012100
2800fdd1
bd38d1f9
4ff0e92d
6843461f
4604b08b
0040f013
4693460d
8050f8dd
9054f8dd
6861d009
0240f021
6a236062
d4fc04d8
90062001
9006e000
04496a21
7969d510
0202f001
b99bb2d3
69607929
0241f3c1
21011d13
f203fa01
0002ea20
e0076160
f0226862
60630340
05426a20
e7e6d5fc
0f00f1b8
44c1d002
0908ea29
0a00f04f
43c8ea4f
97089309
f8cd9707
46d4a014
0f00f1b9
8097f000
0f00f1bc
7baed133
d50507f3
00c4f8d4
2100f440
10c4f8c4
4620465a
f7fe4629
7baafed9
d51007d6
30c4f8d4
2600f423
60c4f8c4
f895792a
4620a000
f3c22103
f3ca0241
f7fe1a01
6920fea8
792e4949
e001f895
f4414001
f3c61300
99090241
3042ea43
90054308
1cdeea4f
f04fe001
786b0c01
0680f003
b912b2f2
0601f108
f647e004
45b176fc
464ebf38
05b39805
0104f040
40d3ea41
ea400ab2
612161c2
07d8796b
ebc644b3
d5120909
9b179a16
92009918
91029301
0040f104
46324639
f8cd4643
19bfc010
ff30f7ff
c010f8dd
f1b8e792
d10c0f03
46139a08
06016a20
6c21d4fc
1b04f843
429818b0
d1f59308
f1b8e782
d10c0f01
46139a07
06086a21
6c20d4fc
0b02f823
429918b1
d1f59307
f1b8e772
f47f0f00
19beaf6f
06016a20
6c22d4fc
2b01f807
d1f742b7
6921e764
52fff421
001ff022
0301f040
7ba96123
d50a07ca
792b7aea
1205f36a
462072ea
f3c34651
f7fe0241
9806fe20
d1062801
f0416861
60620240
04db6a23
b00bd5fc
8ff0e8bd
07c78000
4ff0e92d
f8dd790d
f8dda030
ac099034
0f01f015
4690460e
0890e894
e8bdd103
f7ff4ff0
910abee7
0041f3c5
461a4611
97094623
4ff0e8bd
bd0df7fe
4604b510
f4414613
21104240
fcaef7fe
f4236923
f02050ff
f041011f
61220201
6a03bd10
d406045a
07cb6901
6842d5fc
0340f042
47706043
4ff7e92d
f002784a
b2dd0304
92014604
6842b11d
0710f042
6846e002
0710f026
798b6067
6090f8d4
0507f003
bf0c2d04
2600f446
2600f426
6090f8c4
7a0e790f
0f06f017
f104bf14
f1040094
f0060090
68020302
0cfff003
788fb12b
6207ea42
2580f442
f422e001
7b4b2580
0708f003
b112b2fa
3580f445
f425e001
f0033580
b2fa0720
f445b112
e0015500
5500f425
0710f003
b112b2fa
3500f445
f425e001
f0033500
b2fa0740
f445b112
e0014580
4580f425
0380f003
b117b2df
4200f445
f425e001
89cd4200
13c3f3c5
0743ea42
bf4c07f6
1780f447
1780f427
79086007
f3c0250c
435d0341
0708f104
060cf104
0f00f1bc
8908d003
0287f3c0
788ae000
f8460212
79482025
9025f856
0802f000
f288fa5f
f049b112
e0010a01
0a01f029
a025f846
f89188ca
f3c2b002
7aca0cc7
680cea4f
490bea48
1a92ea4f
c001f891
1b0aea49
9006f891
0808f00c
0a01f109
0208ea4b
0b01f00a
0c4bea42
2025f856
080cea42
8025f846
a009f891
9003f891
c004f891
02c3f3ca
1b19ea4f
7a02ea4f
09c0f3cc
f8919a01
f002c001
f3cc0280
ea4a1800
f00c6a0b
f88d0c03
ea4a2004
ea4c0c0c
f89159c9
ea49c000
f00c4888
ea480903
f3cc1889
b2d20981
1809ea48
1c9cea4f
bf142a00
3220f44f
ea482200
ea4c0c8c
f8470202
f8912025
f01cc00e
bf080f01
c000f891
0070f000
f3ccbf0a
f4421c01
ea427240
2870220c
2025f847
794ad021
1202f3c2
21104620
4240f442
fb90f7fe
f4206920
f02151ff
f043031f
61220201
f0406860
60610120
3025f857
5280f043
2025f847
0025f856
2140f440
1025f846
6861e003
0320f021
46206063
e8bdb003
f7ff4ff0
e92dbec8
460d47f0
7baf7909
6020f89d
f0014604
28060006
469a4690
0941f3c1
0741f3c7
2804d009
2802d00a
200ebf0c
bf0c200a
21002108
201ee004
e0012118
2110201a
23036862
f300fa03
0303ea22
f3c2786a
fa021241
792af000
1200f3c2
4002ea40
60634303
20b0f8d4
fa00200f
ea22f001
7caa0300
00c3f3c2
f101fa00
4620430b
464a2100
30b0f8c4
fc63f7fe
f8d47baa
f01200c4
f1090f01
d0100c02
094cea4f
0308f040
f209fa07
0702ea43
70c4f8c4
00c4f8d4
2100f440
10c4f8c4
ea4fe009
fa07094c
f047f709
ea200108
f8c40701
f1b870c4
d0040f00
46294620
f7ff4652
7babfb6b
d50507da
20c4f8d4
2000f422
00c4f8c4
792b7829
f0014620
f3c30103
f7fe0241
7beafc26
0008f002
b121b2c1
46214628
fb76f7fe
792be004
1240f3c3
60200210
f0037beb
b2ca0180
6862b142
417cf04f
0080f042
f8c46060
e00310b4
f0206860
60610180
0208f003
b918b2d0
f0416821
60220201
792a6920
7100f040
0041f3c2
3140ea41
7b6a6121
0002f002
b119b2c1
f4406960
e0024180
f4206960
61614180
0104f002
b118b2c8
f4416961
e0024000
f4216961
61604000
0f01f012
bf146962
3280f442
3280f422
b10e6162
61e02033
f0017969
2a04020c
6922d103
0180f442
b91ae003
f4206920
61210180
0310f003
b120b2d8
3130f8d4
5280f443
f8d4e003
f4211130
46205280
2130f8c4
f7ff4629
7928fdd7
d50407c3
e8bd4620
f7ff47f0
e8bdbdc4
000087f0
4c0db513
2304480d
22002101
fdd5f003
22002101
f0004620
2101fc37
46202200
fc1cf000
21002301
46209300
460b2250
fc54f000
bf00bd1c
24042000
24041400
47f0e92d
4606460c
4611461d
4620b91a
460b4632
2affe004
4620d106
23004632
47f0e8bd
b9f3f7ff
f0020917
2600090f
ea4f454e
d0234886
21084620
462b2206
fa24f7fe
f4236923
f02050ff
f041011f
61220201
21084620
462b2236
fa16f7fe
21204620
462b4642
fa10f7fe
f4236923
f02050ff
f041011f
61220201
e7d73601
b32f4646
21084620
462b2206
f9fef7fe
f4236923
f02050ff
f041011f
61220201
21084620
462b2239
f9f0f7fe
46204632
462b2120
f9eaf7fe
f4236923
f02050ff
f041011f
61220201
2680f506
e7d83f01
87f0e8bd
47f0e92d
f890461f
7b839004
460d2600
46904604
0941f3c9
03c3f3c3
428b4631
2201d005
f201fa02
31014316
78e0e7f7
010ff000
d1142908
463a4621
f7fe4628
464afbdf
46234682
21354628
f9c6f7fe
230aea40
ea2302b0
ea000200
43322688
290ae015
4620d107
46424629
e8bd464b
f7ff47f0
463abf5b
46214628
fbc0f7fe
ea2000b6
ea060006
ea400688
b2910206
46224628
e8bd463b
f7ff47f0
0000b94e
23004a07
60536013
60d36093
61536113
61d36193
62536213
62d36293
bf004770
46006000
4b04b508
601a2201
ffe8f7ff
20084902
bd086008
460081b4
460081c0
1201eb02
58810112
0100f363
47705081
1201eb02
1002eb00
47706043
1201eb02
1002eb00
b2c86841
eb024770
01111201
f0005840
47700001
7110f501
f850b510
f3634031
f840240b
f8504031
f3623031
f840330d
bd103031
7110f501
3031f850
0208f043
2031f840
f5014770
f8507110
f36f3031
f84003c3
47703031
7110f501
3031f850
0204f043
2031f840
f5014770
f8507110
f36f3031
f8400382
47703031
7110f501
3031f850
0202f043
2031f840
f5014770
f8507110
f0433031
f8400210
47702031
7110f501
3031f850
1304f36f
3031f840
f5014770
f8507110
f36f3031
f8400341
47703031
7110f501
3031f850
0201f043
2031f840
f5014770
f8507110
f36f3031
f8400300
47703031
7110f501
00c1eb00
b2d06842
f5014770
eb007110
684300c1
6042431a
eb024770
01121201
f3635881
50810185
31184770
3021f850
0302f362
3021f840
eb024770
01111201
f0435843
50420202
eb024770
01111201
f36f5843
50430341
eb004770
f5011141
68d85380
000ff362
477060d8
eb003180
60421041
31804770
50420149
eb004770
688b1101
030ff362
4770608b
1141eb00
5080f501
47706082
1141eb00
5080f501
47706102
1141eb00
5380f501
b2806958
eb024770
01111201
f4435843
50427280
eb024770
01111201
f36f5843
50432308
eb024770
01111201
f4435843
50426280
f5014770
f8507112
f0433031
f8400210
47702031
7112f501
3031f850
1304f36f
3031f840
f5014770
f8507112
f0433031
f8400208
47702031
7112f501
3031f850
03c3f36f
3031f840
f5014770
f8507112
f36f3031
f8400341
47703031
7112f501
3031f850
0202f043
2031f840
f5014770
f8507112
f36f3031
f8400300
47703031
7112f501
3031f850
0201f043
2031f840
f5014770
eb007112
684000c1
f5014770
f8507112
f0433031
f8400204
47702031
7112f501
3031f850
0382f36f
3031f840
f5014770
eb007112
604200c1
eb024770
01111201
f36f5843
5043238a
eb024770
01121201
f3635881
50812149
eb024770
01121201
f3635881
508121cb
00004770
21014b03
fa01681a
4302f000
4770601a
41300610
508cf100
5380f500
680a0099
0010f042
47706008
508cf100
5380f500
680a0099
600a2200
00004770
22204b01
4770601a
41300004
508cf100
5280f500
f64f0092
6810733f
ea434003
60111181
f1004770
f500508c
00925280
73fcf64f
40036810
60114319
f1004770
f500508c
00925280
73fbf64f
40036810
0181ea43
47706011
508cf100
5280f500
f64f0092
681073f7
ea434003
601101c1
f1004770
f500508c
00925280
73dff64f
40036810
1141ea43
47706011
21014b03
fa01681a
4302f000
4770601a
2404a008
681a4b02
601a2200
bf004770
2404a008
d1042819
681a4b14
5000f442
281ae021
4b11d104
f4416819
e01a4080
d104281b
68184b0d
4000f440
281ce013
4b0ad104
f442681a
e00c3080
d104281d
68194b06
3000f441
281ee005
4b03d104
f442681a
60182080
bf004770
46008044
d81e280f
f000e8df
08080808
0a0a0a0a
0c0c0c0c
15151515
e0024a0a
e0094b09
68104a09
733ff64f
ea434003
60111181
4b054770
04826818
ea400c90
b28a3181
4770601a
2404a000
2404a004
d81c280f
f000e8df
08080808
0a0a0a0a
0c0c0c0c
13131313
e0024a09
e0074a08
68104a08
73fcf64f
43194003
4a05e006
f64f6810
400343ff
2101ea43
47706011
2404a000
2404a004
d81f280f
f000e8df
08080808
0a0a0a0a
0c0c0c0c
15151515
e0024a0b
e0094a0a
68104a0a
73fbf64f
ea434003
60110181
4a064770
f64f6810
400333ff
2181ea43
6010b288
bf004770
2404a000
2404a004
d81f280f
f000e8df
08080808
0a0a0a0a
0c0c0c0c
15151515
e0024a0b
e0094a0a
68104a0a
73f7f64f
ea434003
601101c1
4a064770
f24f6810
400373ff
21c1ea43
6010b288
bf004770
2404a000
2404a004
d81f280f
f000e8df
08080808
0a0a0a0a
0c0c0c0c
15151515
e0024a0b
e0094a0a
68104a0a
73dff64f
ea434003
60111141
4a064770
f64d6810
400373ff
3141ea43
6010b288
bf004770
2404a000
2404a004
d8072903
00c1eb00
f0437903
71010101
47702000
0001f640
29034770
eb00d807
790300c1
0140f043
20007101
f6404770
47700001
d8072903
00c1eb00
f0437903
71010104
47702000
0001f640
29034770
eb00d807
790300c1
0104f023
20007101
f6404770
47700001
d8072903
00c1eb00
f0437903
71010102
47702000
0001f640
29034770
f840d803
20002031
f6404770
47700001
d8072903
3080f8b0
b29a2001
f001fa00
47704010
47702000
d80d2a03
d80e2902
00c2eb00
0103f001
f0237903
ea420218
710101c1
47702000
0001f640
f6404770
47700003
d80d2a03
d80e2901
00c2eb00
0101f001
f0237903
ea420220
71011141
47702000
0001f640
f6404770
47700002
d8052903
01c1eb00
f3c08888
477000c1
0001f640
eb004770
791a03c1
027ff062
f850711a
47700031
2903b510
4008f89d
2c01d818
f8b0d109
f8a01084
b2d92084
2088f890
1088f880
2c02e00a
f8b0d10a
f8a0108c
b2db208c
2090f890
3090f880
bd102000
0002f640
b082bd10
3081f44f
4770b002
47702014
47702018
47706101
791a6843
0001f042
47707118
791a6843
0001f022
47707118
f0006cc0
47700001
d806291f
22016843
f101fa02
20006299
f2404770
47703001
68986843
68434770
477068d8
4ff0e92d
69406845
b050f8d5
9c096849
0a01f04f
fa00fa0a
ea4a0f96
29010a0b
0907f002
1709f3c2
3883f3c2
6c81f3c2
a050f8c5
3020d101
2900e002
2000bf18
293fb281
8091f200
290068a9
8090f000
0107f002
29023901
f20068ad
f000808d
ea4f0a3f
eb051b0a
f1b8010b
68880f0a
0002f369
68886088
09c0f3c2
00c3f369
68886088
100df367
dd036088
3005f240
8ff0e8bd
f3686888
60883091
f3c26888
f3684882
60884094
f3c26888
f3685842
60885057
f0000e10
f1b80803
d0e50f03
8008f8d1
6901f3c2
6819f369
8008f8c1
080cf010
f1b8d008
d0050f04
0f08f1b8
f1b8d002
d1d10f0c
8008f8d1
689bf36c
8008f8c1
0830f010
f1b8d005
d0020f10
0f20f1b8
f8d1d1c2
f3c28008
f3697901
f010781d
f8c100c0
d0058008
d0032840
d0012880
d1b128c0
f1bc6888
bf180f03
fc0cfa07
709ff366
4463bf18
b1fb6088
f8452e03
d00e300b
0207f002
d0012a04
d1052a06
0420f04a
1404eb05
e002340c
f606fa07
b17c19a4
2000604c
8ff0e8bd
3002f240
8ff0e8bd
3003f240
8ff0e8bd
3006f240
8ff0e8bd
3007f240
8ff0e8bd
2b01684b
6943d102
e0033320
6943b90b
2300e000
2a3fb29a
6840d811
b1816881
f0036882
eb02033f
68811003
f3c16883
f0031209
b9020007
1c50b128
20004770
f2404770
47703002
2b01684b
6943d102
e0033320
6943b90b
2300e000
2a3fb29a
6840d80b
b1516881
f0036882
eb02033f
68811003
0007f001
20004770
f2404770
47703002
68186843
0001f000
68434770
f3c06818
47701003
460db538
0103f010
d1104604
f00b2218
68aafac5
6869682b
f4226023
f020707f
42930303
60a26061
608bd103
2000e001
4620bd38
291fbd38
6843d80a
fa226a9a
f011f101
f64f0f01
bf1870ff
e0012000
3001f240
4770b200
2b1fb28b
6843d808
695a2001
f101fa00
61594311
47702000
3001f240
00004770
b570291f
6840d83a
2c006884
2b00d036
f5b2d034
d8316f80
010eb382
eb036884
3b041302
4b1751a3
eb044298
d1020506
0320f041
4b14e004
d1054298
0310f041
1403eb04
606c340c
23002402
739ff364
731df364
639bf364
6319f364
3391f364
00929c04
0302f364
f3623a01
60ab130d
fa032301
6341f101
bd702000
3005f240
bf00bd70
44030000
24078000
2b1fb28b
6843d80a
f8d32001
fa002800
4311f101
1800f8c3
47702000
3001f240
b5304770
b0856903
2b004604
8162f000
f8d16841
07e95800
2100d507
ffe0f7ff
46206923
22004669
07aa4798
2101d508
f7ff4620
6923ffd5
46694620
47982201
d508076b
46202102
ffcaf7ff
46206923
22024669
07284798
2103d508
f7ff4620
6923ffbf
46694620
47982203
d50806e9
46202104
ffb4f7ff
46206923
22044669
06aa4798
2105d508
f7ff4620
6923ffa9
46694620
47982205
d508066b
46202106
ff9ef7ff
46206923
22064669
06284798
2107d508
f7ff4620
6923ff93
46694620
47982207
d50805e9
46202108
ff88f7ff
46206923
22084669
05aa4798
2109d508
f7ff4620
6923ff7d
46694620
47982209
d508056b
4620210a
ff72f7ff
46206923
220a4669
05284798
210bd508
f7ff4620
6923ff67
46694620
4798220b
d50804e9
4620210c
ff5cf7ff
46206923
220c4669
04aa4798
210dd508
f7ff4620
6923ff51
46694620
4798220d
d508046b
4620210e
ff46f7ff
46206923
220e4669
04284798
210fd508
f7ff4620
6923ff3b
46694620
4798220f
d50803e9
46202110
ff30f7ff
46206923
22104669
03aa4798
2111d508
f7ff4620
6923ff25
46694620
47982211
d508036b
46202112
ff1af7ff
46206923
22124669
03284798
2113d508
f7ff4620
6923ff0f
46694620
47982213
d50802e9
46202114
ff04f7ff
46206923
22144669
02aa4798
2115d508
f7ff4620
6923fef9
46694620
47982215
d508026b
46202116
feeef7ff
46206923
22164669
02284798
2117d508
f7ff4620
6923fee3
46694620
47982217
d50801e9
46202118
fed8f7ff
46206923
22184669
01aa4798
2119d508
f7ff4620
6923fecd
46694620
47982219
d508016b
4620211a
fec2f7ff
46206923
221a4669
01284798
211bd508
f7ff4620
6923feb7
46694620
4798221b
d50800e9
4620211c
feacf7ff
46206923
221c4669
00aa4798
211dd508
f7ff4620
6923fea1
46694620
4798221d
d508006b
4620211e
fe96f7ff
46206923
221e4669
2d004798
211fda08
f7ff4620
6923fe8b
46694620
4798221f
bd30b005
2a1f69ca
6142b530
2401d86e
fa046843
4c38f202
42a364da
4c37d104
432a6825
e0086022
42a34c35
f8b3d105
4322482a
f8a3b292
684a282a
d1032a01
fa026944
631af204
2a01688a
6944d103
f204fa02
68ca619a
d1082a01
2a1f8a82
f893d805
f0422828
f8830201
690a2828
d1032a01
fa026944
621af204
2a01680a
6940d103
f200fa02
694b639a
d1302b01
1e486989
d82c2806
f000e8df
130e0904
00221d18
68194b17
0101f041
4b15e01c
f042681a
e0170102
68184b12
0108f040
4b10e012
f0416819
e00d0110
681a4b0d
0120f042
4b0be008
f0406818
e0030140
681a4b08
0180f042
e0026019
3001f240
2000bd30
bf00bd30
44030000
4611000c
24078000
46008058
4801b082
4770b002
02000001
f44f2220
e8806c80
47701004
d806291f
22016843
f101fa02
200062d9
f2404770
47703001
4604b538
6941460d
fde4f7ff
69614620
ffeaf7ff
791a6863
0001f022
69627118
d8172a1f
b91968a9
fa002001
61d8f002
b9196869
fa002001
6358f002
b9196829
fa002001
63d8f002
b9196929
fa002001
6258f002
fa012101
64daf202
6843bd38
f8d32001
fa002800
4010f001
694b4770
b5702b07
68ccd819
d1082c01
f5026842
009e5284
fa0468d5
432cf406
690960d4
d10d2901
f5006840
009b5284
330368d0
f103fa01
60d14301
f240e002
bd702001
bd702000
f5036843
20015384
fa00695a
430af101
2000615a
20244770
00004770
2b07694b
6203b5f0
680ed860
d85d2e03
f5046844
692a5584
b2d2401a
d0582a01
eb006880
ea4f2003
8a870cc3
0238f00c
073ff027
8282433a
f4278a87
f442627c
82877700
f0067e02
f0220603
43160203
68ca7606
d1052a01
009e68e8
f206fa02
60ea4302
28016908
f504d108
009e5284
360368d5
f006fa00
60d04328
25014a17
fa056810
4303f303
f5046013
684c5384
2c01689d
6888d120
2801694a
689cd10e
0108f102
fa003210
fa00f101
ea24f002
ea650101
40080000
e00d6098
32086899
f402fa04
0404ea21
e005609c
200af240
f240bdf0
bdf0200b
bdf02000
46110004
d80a2903
f001e8df
08060402
47706102
47706142
47706182
477061c2
b912b570
220af240
7b8de0e2
1401f3c5
d0f72c03
0581f3c5
d0f32d03
8990898e
000bf366
7b488190
0030f010
2810d006
2820d004
2830d002
80bff040
7b507b4e
1601f3c6
1005f366
7b487350
00c0f010
2880d006
2840d004
28c0d002
80b0f040
7b507b4e
f36609b6
73501087
7b907b8e
0000f366
7b8e7390
f3c6b2c0
f3660640
73900041
f0107b88
d003000c
d0012804
d1b72808
f3657b90
73900083
f0107b88
d0030030
d0012810
d1ab2820
f3647b90
73901005
b2c07b8c
1480f3c4
1086f364
7b8c7390
09e4b2c0
10c7f364
7bcc7390
f3647bd0
73d00000
b2c07bcc
0440f3c4
0041f364
7bcc73d0
f3c4b2c0
f3640480
73d00082
b2c07bcc
04c0f3c4
00c3f364
7bcc73d0
f3c4b2c0
f3641400
73d01004
b2c07bcc
1440f3c4
1045f364
7bcc73d0
f3c4b2c0
f3641480
73d01086
7c107c0c
0002f364
7c4c7410
f3c47c50
f3640445
74500046
8a108a0c
04c5f3c4
00c8f364
690c8210
34c5f3c4
f73f2c2f
6910af53
30d4f364
8a4c6110
1445f3c4
f73f2c2f
8a50af49
104af364
7ccc8250
f3c47cd0
f36404c2
74d000c5
b2c07ccc
1480f3c4
1086f364
7ccc74d0
09e4b2c0
10c7f364
684874d0
6889b178
b1796050
b1136091
2200601a
6013e00c
f44fe7fb
e0077202
2202f240
f44fe004
e0017201
2205f240
bd70b210
2b07694b
d819b570
2c01684c
6842d109
5284f502
68d5009e
fa043601
432cf406
688c60d4
d1092c01
f5056845
009b5284
330268d5
f403fa04
60d4432c
4070e8bd
be45f7ff
d8082907
f5036843
69025084
fa002001
4010f001
f2404770
47702001
460db538
0103f010
d10c4604
f00a2224
682bfe2d
68a96868
606068ea
60a16023
462060e2
2000bd38
2907bd38
6843d80a
5384f503
691a2001
f101fa00
61194311
47702000
2001f240
29074770
f200b570
688480e9
eb048995
68d82301
000bf365
7b5360d8
0030f013
2810d006
2820d004
2830d002
80caf040
2001eb04
68c57b56
1601f3c6
350df366
03c0f013
d00660c5
d0042b80
d0022b40
f0402bc0
eb0480ba
7b552301
09ad68d8
308ff365
68d860d8
f3657b95
60d84010
68d87b95
0540f3c5
4051f365
7b9360d8
0030f013
2810d006
2820d004
f240d002
bd70200a
2001eb04
1601f3c3
f01368c5
f366030c
60c55515
2b04d003
2b08d001
0209d1ed
f1001860
7b960308
f3c6685d
f3660681
605d4593
685d7b96
1680f3c6
5596f366
7b96605d
09f6685d
55d7f366
685d605d
f3667bd6
605d6518
685d7bd6
0640f3c6
6559f366
7bd6605d
f3c6685d
f3660680
605d659a
685d7bd6
06c0f3c6
65dbf366
7bd6605d
f3c6685d
f3661600
605d751c
685d7bd6
1640f3c6
755df366
7bd6605d
f3c6685d
f3661680
605d759e
69037c15
0302f365
7c556103
f3c56903
f3650545
6103234e
69038a15
05c5f3c5
03c8f365
69156103
35c5f3c5
dc8e2d2f
f3656903
610333d4
f3c58a55
2d2f1545
6903dc85
535af365
7cd56103
f3c56903
f36505c2
610363dd
69037cd5
1580f3c5
739ef365
7cd56103
09ed6903
73dff365
68536103
6043b163
b1636893
50626083
bd702000
7002f44f
f240bd70
bd702002
7001f44f
f240bd70
bd702005
2001f240
b570bd70
f5036843
46045184
6a0168cd
1cda008b
f202fa25
f303fa25
07d3431a
f7ffd51c
2100fd33
f7ff4620
6a22fd0c
fa250090
07c9f100
69a3d504
4620b113
47982100
00906a22
fa251cc1
07dbf301
69e3d504
4620b113
47982100
00906a22
fa251c41
07d8f301
6866d50d
5384f506
68d82601
f101fa06
60d94301
b1136963
21004620
6a224798
1c810090
f501fa25
d50d07eb
f5056865
25015384
fa0568d8
4301f101
692360d9
4620b113
47982100
b082bd70
3081f44f
4770b002
20002308
0003f363
f3612102
22401005
108cf362
f3632304
4770304f
2b07694b
684ad816
d1062a01
f5016841
009b5084
1c5868c1
688ae008
d10c2a01
f5016841
009b5084
1c9868c1
f000fa02
47704008
2001f240
20004770
694b4770
d8152b07
2a0168ca
6841d105
5084f501
009868c1
690ae008
d1092a01
f5016841
009b5084
1cd868c1
f000fa02
47704008
47702000
b5f02a07
4b15d824
681d2401
f402fa04
601c432c
684d6844
5384f504
68982d01
689ed108
0708f102
fa054306
ea66f507
609d0505
29016889
f504d10d
32105384
fa01689c
4320f102
0201ea60
e002609a
2001f240
2000bdf0
bf00bdf0
46110004
f64f4b04
801a72ff
068b6d81
2000d5fc
bf004770
46188068
b390b538
f8d44c1a
f0455080
f8c40580
4c185080
15fff240
b1f18025
1014f8bd
4915008c
5c40f831
052c800c
501cf8bd
0ce40252
03c3ea42
3445ea44
4c40f821
3c04f821
1010f8bd
3018f8bd
f042018a
f0030208
430a013f
f243e001
4b0712c1
f7ff801a
2000ffc1
2001bd38
bf00bd38
24048400
46188068
46188048
46188040
b920b570
f5b1b119
f2407f96
4b428082
f1f3fbb1
fbb22901
d90ef2f3
d90e2903
d90e2907
d90e290f
d90e291f
d90e293f
bf8c297e
23012300
2307e00a
2306e008
2305e006
2304e004
2303e002
2302e000
fa052501
4d31f603
f403fa01
f8d51e73
f0466080
f8c50680
4d2d6080
16fff240
b2a429c8
802eb29b
f011d907
f1a50101
bf180520
4100f44f
2cfa8029
d9104925
0535880e
3a010cee
00d24d23
2343ea42
43350864
878b800d
018a1e61
040af042
f1a4e029
2e3106c9
880ed811
0cee0535
3a014d19
800d4335
00d10864
ea414a17
1e612343
018b8013
0408f043
4d14e013
802e2600
052d880d
0595ea6f
ea6f3a01
800d4555
00d13c01
ea414a0c
01a12343
f0418013
4b0b0409
f7ff801c
2000ff2d
2001bd70
bf00bd70
000f4240
24048400
46188068
46188008
ffffa000
46188044
46188048
46188040
f2404b02
801a12ff
47702000
46188068
f2434b02
801a12f9
47702000
46188040
f2434b02
801a12c9
47702000
46188040
881a4b04
5093f442
0114f040
20008019
bf004770
461880c0
f2414b02
801a2244
47702000
461880c0
4b05b140
72fff64f
6d81801a
d5fc06ca
47702000
47702001
461880e8
b1f0b538
f2404c10
802515ff
f8bdb1a9
02c95010
ea41005b
01ad2202
430ab2d9
0504f045
5c28f824
2c24f824
2014f8bd
3c284b06
34040091
f7ff8019
2000ffd3
2001bd38
bf00bd38
461880e8
461880c8
47f0e92d
4691460e
28004607
809bf000
429a4b4e
484ed00a
d0074282
4a4e494d
45a94d4e
4614bf14
e000460c
46304c49
ffe2f009
484a4601
f8eaf00a
f00a4605
f009f9f9
4601ffdd
f0094628
2100ff23
f9bef00a
4628b130
fa12f00a
a10cf8df
e004b286
fbb34b3f
b2b6f6f6
4650469a
ffc2f009
46204605
ffbef009
46284601
f8c6f00a
f9f4fbb9
f00a4604
fa1ff9d3
4620f880
fc74f009
46404604
f009460d
4602fc5d
4620460b
f0094629
2200fb09
f0094b2d
f009fcb9
492cfec9
b280458a
3001d101
f5b6b280
d3047f90
1e5e0933
2304b2b6
f1a6e019
2a300260
08f1d804
b2961e4a
e0102303
d00c2e48
0324f1a6
d8042b0c
1e4a0871
2301b296
3e01e005
2300b2b6
2302e001
4a192611
ea4f021b
f2400e49
801111ff
1c88ea4f
26c6ea43
f98efa5f
f04c4913
00800804
0609ea46
8c28f822
6c24f822
46388008
ff2af7ff
e8bd2000
200187f0
87f0e8bd
00927c00
0124f800
000ea600
000f4240
0249f000
4c8ca000
04099800
40d00000
04650000
461880e8
461880c8
f2404b02
801a12ff
47702000
461880e8
f2434b02
801a12f9
47702000
46188080
f2434b02
801a12c9
47702000
46188080
f2404b02
801a12ff
47702000
461880a8
4b05b140
72fff64f
6d81801a
d5fc0709
47702000
47702001
461880a8
b368b538
f2404c17
802515ff
f8bdb301
49154014
f83100a5
800d4c80
b2ac0065
501cf8bd
f4240252
ea4254e0
ea4403c3
f8212485
f8214c80
f8bd3c04
f8bd1010
018a3018
0208f042
013ff003
e001430a
12c1f243
801a4b05
ffc4f7ff
bd382000
bd382001
461880a8
46188088
46188080
b918b570
f5b1b111
d97e7f96
4b414e40
f1f6fbb1
14fff240
801c2901
f2f6fbb2
2903d90e
2907d90e
290fd90e
291fd90e
293fd90e
297ed90e
2600bf8c
e00a2601
e0082607
e0062606
e0042605
e0022604
e0002603
fa012602
b2acf506
fa052501
1e5ef306
b2b329c8
4029d905
bf184d2a
4100f44f
2cfa8029
d9134928
f24e880e
007635fe
00d23a01
ea424035
08642343
55a0f445
f8a1800d
1e61307c
f042018a
e02c040a
06c9f1a4
d8132e31
f24e880e
007635fe
3a014035
55a0f445
0864800d
4a1700d1
2343ea41
80131e61
f043018b
e0140408
26004d10
880e802e
35fef24e
40350076
f4453a01
800d5580
00d13c01
ea414a0b
01a12343
f0418013
4b090409
f7ff801c
2000ff37
2001bd70
bf00bd70
000f4240
461880a8
46188088
46188008
46188084
46188080
6001b110
47702000
47702001
6041b110
47702000
47702001
6081b110
47702000
47702001
60c1b110
47702000
47702001
6101b110
47702000
47702001
6141b110
47702000
47702001
6c43b128
0101ea23
20006441
20014770
b0824770
93012300
d8182903
f001e8df
0e0a0602
f0136d83
e00a0f20
f0126d82
e0060f08
f0116d81
e0020f10
f0106d80
d0010f40
e0012000
7001f241
98019001
4770b002
6c43b120
64414319
47702000
47702001
4615b538
b9084604
d93e2a3f
68d84b20
bf480782
2905086d
e8dfd837
3603f001
241b1207
f36f6aa3
e0240303
21004620
ffbdf7ff
f241b110
bd387001
20026aa3
4620e017
f7ff2103
2800ffb2
6aa3d1f3
e00e2003
21014620
ffa9f7ff
d1ea2800
20046aa3
490be005
07536a4a
6aa3d5e3
f3602005
62a30303
05c86da1
6aa2d5fc
1209f365
200062a2
2001bd38
bf00bd38
24048600
24041400
b929b178
60432302
f4416c41
e0067200
d1082901
60432308
f4416c41
64426200
2001e001
20004770
b1884770
7380f04f
60c3b921
f3616c43
e0065355
6180f04f
61016083
f4426c42
64431300
47702000
47702001
b939b188
f44f6c42
f36143c0
64424292
e00660c3
4360f44f
6c416083
4192f36f
20006441
20014770
b1284770
f3616a83
62831309
47702000
47702001
b1c8b510
6981b121
7100f441
e0036181
f3616984
61842449
69c2b122
5180f042
e00361c1
f36269c1
61c1711c
f3636982
618202c8
bd102000
bd102001
6a83b128
5319f361
20006283
20014770
b1284770
f3616983
618323ce
47702000
47702001
69c3b128
631bf361
200061c3
20014770
b1284770
f3616a83
628323d0
47702000
47702001
6c03b168
f443b111
e0017300
2349f361
6c016403
0105f362
20006401
20014770
b1f04770
b122b969
f04269c2
61c15100
69c1e003
715df362
69c261c1
02c6f363
b122e00c
f04269c2
61c14180
69c1e003
719ef362
69c261c1
228df363
200061c2
20014770
00004770
2903b908
2903d929
e8dfd827
0b02f001
4b131813
f4416a19
621a3280
f36f6a41
e0145156
6a194b0e
2280f441
6a41621a
e0012201
22026a41
5156f362
4b08e007
f4426a1a
62193100
f4436a43
624101c0
02996d83
2000d5fc
20014770
bf004770
24048100
4604b510
2c002001
69a3d038
62e0f043
60a061a2
d82d2904
f001e8df
180d0a03
f04f0021
61236380
f36f69a0
e020601a
210169a0
4620e01b
f7ff2100
b110fe7c
7001f241
69a0bd10
e0102102
21034620
fe71f7ff
d1f32800
210369a0
4620e007
f7ff2101
2800fe68
69a0d1ea
f3612104
61a0601a
04d06da2
2000d5fc
0000bd10
5380f44f
b5702901
460d4604
61434616
d302d019
d1232902
2103e010
fe4bf7ff
f241b110
bd707001
880a490e
f043b293
800a0240
f3606aa1
e007715e
f7ff2103
2800fe3a
6aa1d1ed
715ef365
6fe062a1
5380f44f
00c4f366
612367e0
bd702000
bd702001
4113801c
d0402800
d83e290b
f001e8df
100c0906
1f1c1a17
37302a24
7300f44f
f04fe02b
e0285300
6280f04f
e0046002
6300f44f
f44f6083
61025200
f44fe023
e01a5300
e00b2140
2180f44f
f04fe008
61026280
e0032108
6380f04f
21016103
e0106081
1100f44f
f44f6081
e7e43280
6280f04f
f44f6102
60031300
6a03e003
2180f443
20006201
20014770
28004770
290dd047
e8dfd845
0f07f001
20191512
2f2c2a27
3e3a3431
7280f04f
6c4360c2
1100f443
e0326441
7100f44f
f04fe029
e0265100
6380f04f
e00b6043
f4436c43
64412180
41c0f44f
f44fe011
60c26200
43c0f44f
e01a6143
5100f44f
2140e011
f44fe005
e0022180
e0002108
60c12101
f44fe00d
60c21200
3380f44f
f44fe7ea
60411100
6a03e003
4392f36f
20006203
20014770
00004770
4b04b908
2801e002
4b03d0fb
f3c08818
47703080
46188070
461880f0
881a4b05
bf0c2801
0208f042
0208f022
2000801a
bf004770
46188040
881a4b05
bf0c2801
0204f042
0204f022
2000801a
bf004770
46188040
881a4b05
bf0c2801
0210f042
0210f022
2000801a
bf004770
46188040
881a4b05
bf0c2801
0208f042
0208f022
2000801a
bf004770
461880c0
881a4b05
bf0c2801
0204f042
0204f022
2000801a
bf004770
461880c0
881a4b05
bf0c2801
0210f042
0210f022
2000801a
bf004770
461880c0
881a4b05
bf0c2801
0208f042
0208f022
2000801a
bf004770
46188080
881a4b05
bf0c2801
0210f042
0210f022
2000801a
bf004770
46188080
881a4b05
bf0c2801
0204f042
0204f022
2000801a
bf004770
46188080
b959b1d8
b9222102
6c436041
2349f362
6001e011
f4426c42
e00c7300
d10e2901
b9222308
6c436043
23cbf362
6003e003
f4416c41
64436300
2001e001
20004770
e92d4770
9e0943f8
8020f89d
46174689
4604461d
2e0fb910
80adf240
46294620
fd4cf7ff
0f04f1b8
80a5f200
f008e8df
35175003
b93d006a
f36569e0
61e00002
054a6da1
e069d5fc
f0402d01
69e0808c
10c9f36f
6da161e0
d5fc050b
4620e077
f7ff2103
b118fcb6
7001f241
83f8e8bd
69e0b945
f3622202
61e00002
05486da1
e04bd5fc
d16e2d01
210269e0
10c9f361
6da361e0
d5fc0519
4620e059
f7ff2101
2800fc98
b945d1e0
230369e1
0102f363
6da261e1
d5fc0552
2d01e030
69e3d153
f3622203
61e313c9
05036da0
e03ed5fc
21004620
fc7df7ff
d1c52800
69e1b945
f3622201
61e10102
05586da3
e015d5fc
d1382d01
f36569e3
61e313c9
05016da0
e024d5fc
69e3b9b5
f3622204
f04f0302
61e36080
6da16120
d5fc054a
f36669e2
61e202c6
b11769e3
735df36f
f043e01a
e0175300
d1162d01
220469e3
13c9f362
6080f04f
612061e3
050b6da1
69e2d5fc
228df366
69e361e2
f36fb117
e001739e
4380f043
462061e3
464a4629
ff28f7ff
e8bd2000
200183f8
83f8e8bd
f44fb1c8
b94163c0
6c4360c3
33cff361
6c426443
4210f361
f04fe00a
60836180
6c426101
4300f442
6c416443
3280f441
20006442
20014770
b5704770
461e460d
b9084604
d92d2b0f
5380f04f
60e32a01
d10a4620
f7ff4611
b110fbfe
7001f241
69a1bd70
4192f360
2100e007
fbf3f7ff
d1f32800
f44069a0
61a12180
03516da2
69a3d5fc
43d6f366
69a061a3
f440b115
e0010000
50d7f365
5180f04f
60a161a0
bd702000
bd702001
d8382804
28033801
e8dfd82e
0d02f000
4b1a2318
21036a18
0002f361
6a1a6218
0008f042
e01f6218
6a5a4b14
f3612104
625a0202
f0406a58
625a0208
4b0fe014
21056a98
0002f361
6a9a6298
0008f042
e0096298
6ada4b09
f3612106
62da0202
f0406ad8
62da0208
69594b05
0201f041
2000615a
20014770
bf004770
24048600
24048000
2903b180
6e83d80e
0342f361
6e816683
0201f041
6e836682
d5fc031b
f3c06e80
477000cf
47702001
b1a0b510
2480b93a
3300f44f
6084b109
60c4e007
f44fe009
f44f7280
b1192380
61036082
bd102000
614360c2
2001e7fa
b160bd10
60c32308
b2c96a02
0207f361
6180f04f
61016202
20006083
20014770
00004770
460fb5f8
461e4615
b9104604
d8072b3f
6c43e029
41c0f44f
2080f443
60e16460
681a4b13
0000f442
b9456018
21024620
fb3df7ff
6aa2b9c8
228af365
f04fe005
61216180
f4436aa3
62a26280
03826da0
6aa1d5fc
21d0f366
462062a1
f7ff4639
2000fbc5
2001bdf8
f241bdf8
bdf87001
46008044
4615b538
b9104604
d8042a0f
f04fe02b
60436380
48166143
29016802
3380f422
d00e6003
2902d306
6801d11d
3280f441
e00e6002
6080f04f
6a616120
71dff36f
4620e006
faf9f7ff
6a63b978
4100f043
69e26261
6080f04f
621bf365
602061e2
20006120
2001bd38
f241bd38
bd387001
46008014
4615b538
b9104604
d8032a3f
f44fe034
60437300
d82f2903
f001e8df
1a110602
f36f6aa1
e01a4153
21014620
facbf7ff
f241b110
bd387001
22016aa1
4620e00d
f7ff2100
2800fac0
6aa1d1f3
e0042202
6080f04f
6aa16120
f3622203
62a14153
04196da3
6aa0d5fc
7100f44f
5019f365
602162a0
bd382000
bd382001
460db570
4604461e
2b3fb910
e042d803
5300f04f
2a036043
e8dfd83d
0e02f002
46202017
f7ff2100
b110fa90
7001f241
6c21bd70
1188f360
4620e018
f7ff2103
2800fa84
6c21d1f2
e00d2201
21014620
fa7bf7ff
d1e92800
22026c21
f04fe004
61206080
22036c21
1188f362
6da36421
d5fc0458
f3666c20
64200005
b1156c21
7100f441
f365e001
f04f2149
64215200
60222000
2001bd70
b570bd70
461d460e
b9104604
d8072b0f
f04fe04c
60c37380
f4406c40
64611100
d8432a05
f002e8df
1b120703
69a32d24
33d1f36f
4620e02c
f7ff2100
b110fa3a
7001f241
69a3bd70
e01f2001
21034620
fa2ff7ff
d1f32800
200269a3
4620e016
f7ff2101
2800fa26
69a3d1ea
e00d2003
21034620
fa1df7ff
d1e12800
200469a3
f04fe004
61226280
200569a3
33d1f360
6da161a3
d5fc048b
f36569a2
61a222ce
46314620
fa8ff7ff
bd702000
bd702001
9f06b5f8
461d4616
b9104604
d8062f3f
f44fe052
60c36300
40c0f44f
29046160
e8dfd84a
0703f001
00271b12
f36f69a3
e01d0302
21034620
f9e3f7ff
f241b110
bdf87001
220269a3
4620e010
f7ff2101
2800f9d8
69a3d1f3
e0072201
21004620
f9cff7ff
d1ea2800
220369a3
0302f362
e00261a3
4180f44f
6da06121
d5fc0582
f36769a1
61a101c8
b11669a3
7300f443
f366e001
61a32349
b11569e2
5280f042
f365e001
f44f721c
f44f6000
61e25100
612160a0
bdf82000
bdf82001
4788b508
0000bd08
460bb508
28064611
e8dfd852
1004f000
3a2f241c
4a270045
02406a10
6a10d403
0080f440
2b006210
200ad142
4a21e03e
02806a10
6a10d4f7
1080f440
6a106210
1000f440
4a1be7ee
02c06a10
6a10d4eb
1080f440
4a17e7e6
03006a10
6a10d403
2000f440
bb1b6210
e01f2002
6a104a11
d4030340
f4406a10
62102080
480eb9c3
4a0ce014
03806a10
6a10d403
3000f440
b96b6210
e00920fa
6a104a06
d40303c0
f4406a10
62103080
2096b913
ffa4f7ff
bd082000
24048100
002625a0
4604b510
2a3fb920
290fd806
e091d804
f36f6a03
62034392
f3626a20
62203011
f200290d
e8df8087
0a07f001
2e261e0d
4f463e36
756a6158
22016a23
6a23e067
e0642202
21034620
f91bf7ff
f241b110
bd107001
88014838
f043b28b
80020240
22036a23
2200e053
21012002
ff6af7ff
22046a23
2001e04b
46012200
ff62f7ff
22056a23
2200e043
21012006
ff5af7ff
22076a23
2200e03b
21012004
ff52f7ff
22086a23
2200e033
21012005
ff4af7ff
22096a23
4620e02b
f7ff2101
2800f8e2
6a23d1c5
e022220a
21034620
f8d9f7ff
d1bc2800
220b6a23
4620e019
f7ff2103
2800f8d0
6a23d1b3
e010220c
21004620
f8c7f7ff
d1aa2800
220d6a23
4620e007
f7ff2102
2800f8be
6a23d1a1
f362220e
e008230b
21034620
f8b3f7ff
d1962800
f4416a21
62236370
f4406a20
62212180
bd102000
bd102001
4113801c
4604b510
d02f2800
29043902
e8dfd82c
0703f001
001b120b
20024b14
e01b69da
20034b12
e01769da
21404b11
4b0f8019
69da2004
2200e010
21012002
fee4f7ff
20054b0a
e00769da
22002001
f7ff4601
4b06fedb
200669da
0202f360
6da261da
dafc2a00
bd102000
bd102001
24048100
4113801c
47706101
47706141
47706501
477064c1
47706201
47706241
47706281
477062c1
43196bc3
013ff001
477063c1
f0036bc3
ea22023f
63c10101
64c14770
65014770
04094770
47706541
65810409
65414770
65814770
66814770
66c14770
00004770
60d84b01
bf004770
24048400
60984b01
bf004770
24048400
64984b01
bf004770
24048400
64584b01
bf004770
24048400
43196803
47706001
ea236803
60010101
47702000
200060c1
69034770
0304f361
20006103
69034770
4314f361
20006103
6a034770
62014319
47702000
ea236a03
62010101
47702000
47706a00
47706b80
200063c1
69434770
0305f361
20006143
69434770
230bf361
20006143
69434770
330ff361
20006143
69434770
6319f361
20006143
69434770
5315f361
20006143
69434770
639bf361
20006143
69434770
43d3f361
20006143
69434770
5397f361
20006143
68434770
0300f361
20006043
68434770
0342f361
20006043
68434770
0342f361
20006043
00004770
f44f4b02
669a3200
bf004770
24048400
f2002815
e8df80cf
0016f010
00290022
00370030
004a003e
00580051
00700060
00780068
00890080
009b0092
00ad00a4
00bb00b6
495c00c4
60082001
6a42485b
0301f042
68016243
5200f041
4857e0a9
f0426882
60810101
e01a2302
68814853
0302f041
23046083
4850e013
f0436883
60820204
e00c2308
6882484c
0108f042
23106081
4849e005
f0436883
60810110
4a452320
68036013
1280f443
4b43e081
f4416819
601a1200
e0352240
680a493f
1000f442
22806008
493ce02e
f4406808
600b1300
7280f44f
4838e026
f4436803
60021200
7200f44f
4b34e01e
f4416819
60180080
6280f44f
4b30e016
f442681a
60191100
6200f44f
492ce00e
f4406808
600a1200
5280f44f
4828e006
f0426802
60037300
5200f44f
e0424823
f44f4b22
60184080
68014821
2280f441
491ee039
4000f44f
481d6008
f4426802
e0303280
481a4a19
3180f44f
68036011
6280f043
4815e027
3200f44f
48146002
f0436803
e01e6200
f44f4b10
60182080
6801480f
5280f041
480de015
f0426802
e0107280
f44f4b09
60184000
68014808
3200f441
4b05e007
f44f4805
601a4200
f4416801
60022200
47702000
12080004
24048100
699a4b07
0284f360
7080f5a3
6a03619a
0302f361
6a016203
d5fc070a
bf004770
24048100
68184b01
bf004770
1208000c
2300b082
28159301
e8dfd866
0d0bf000
1513110f
27211c17
423b2d34
504a5e45
5e5e6556
e0212001
e0372002
e0352004
e0332008
e0312010
e02f2020
22104927
204063ca
4b25e02a
63d82020
e0252080
22404922
f44f63ca
e01f7080
20804b1f
f44f63d8
e0197000
6080f44f
491b4a1c
63c86010
4919e030
7280f44f
f44f63ca
e00b6000
f44f4b15
63d97100
5080f44f
f44fe004
e0015000
4080f44f
60184b10
490fe01a
3080f44f
21086008
4b0ce00a
3200f44f
2104601a
4809e004
2280f44f
21026002
63d14a05
4b05e006
f44f4903
60184000
92016b8a
4770b002
24048100
12080008
f2002815
e8df80ac
170bf000
1f1d1b19
3d352e27
5d55454d
81786f66
a198938a
20014950
48506008
f36f6a42
62420200
f36f6801
e091715d
e0062202
e0042204
e0022208
e0002210
4b462220
601a4846
f36f6801
e0815114
68014843
5155f36f
21406001
4b40e035
f36f681a
601a5255
e02e2180
6801483c
5155f36f
f44f6001
e0267180
681a4b38
5255f36f
f44f601a
e01e7100
681a4b34
5296f36f
f44f601a
e0166180
68014830
5155f36f
f44f6001
e00e6100
6801482c
5155f36f
f44f6001
e0065180
681a4b28
6259f36f
f44f601a
48245100
4923e042
4080f44f
48226008
f36f6801
e0394192
481f4b1e
4200f44f
6801601a
4110f36f
491ae030
3080f44f
48196008
f36f6801
e027619a
48164b15
3200f44f
6801601a
61dbf36f
4911e01e
2080f44f
48106008
f36f6801
e015711c
6801480d
6118f36f
4b0ae010
f44f480a
601a4200
f36f6801
e0074151
48064b05
4200f44f
6801601a
41d3f36f
20006001
bf004770
12080000
24048100
681a4b02
60184310
47702000
24048100
681a4b03
0000ea22
20006018
bf004770
24048100
4605b538
481f460c
3100f44f
fd3bf7ff
695a4b1d
6040f042
69596158
7240f041
6958615a
0140f440
695a6159
1040f442
69596158
2200f441
6958615a
300ff365
695d6158
250bf364
6c1c615d
44d3f36f
6859641c
0100f36f
4b0c6059
f012681a
461c0508
4807d1f9
f7ff213f
4806fcf7
f3656841
60410142
f0136823
d1fb0004
bf00bd38
24048400
24048100
1208001c
2600b5f7
4e389601
402cf89d
5030f89d
60372706
68774e35
0742f360
98016077
48331c46
68069601
d5f80770
6946482f
669bf361
69416146
6119f362
69426141
5297f363
69436142
1020f89d
5315f361
69436143
2024f89d
43d3f362
69416143
4110f365
2d016141
d1076943
3200f443
68416142
4110f36f
e0026041
4351f364
481a6143
69432c01
f443d10e
61413100
f36f6843
60434310
6c04b97d
2034f89d
44d3f362
e0086404
4351f364
68446143
2028f89d
4410f362
4c0c6044
f0406960
6161013f
213f480b
fc7af7ff
f0436863
60620201
4b069801
91011c41
0711681a
2000d5f8
bf00bdfe
24041424
24048100
1208001c
24048400
4803b508
3100f44f
fc7bf7ff
bd082000
24048400
2901b190
6a41d10b
615ef362
6a826241
721cf363
4300f04f
60036282
f04fe002
60434300
47702000
47702001
6803b120
60014319
47702000
47702001
6803b128
0101ea23
20006001
20014770
b9084770
d9122aff
30a4f8d0
f443b111
e0017380
2308f361
30a4f8c0
10a4f8d0
f362b2d2
f8c00107
200010a4
20014770
28004770
818ef000
f200290b
e8df818b
000cf011
00420027
0096007b
00e800c1
015b00ed
012400f2
2a010184
d10b6983
0201f043
68036182
0120f043
f8d06001
f04220a0
e05c0201
0300f36f
68016183
1145f36f
f8d06001
f36f20a0
e0500200
68032a01
f443d10c
60024280
f4436803
60011180
f4426802
60032300
47702000
43d3f36f
68016003
318ef36f
68036001
5314f36f
2a01e7f1
d1196b43
0101f043
f8d06341
f44220a0
f8c05380
f8d030a0
f44110a0
f8c06200
f8d020a0
f44330a0
f8c04100
f8d010a0
f44220a0
e0184280
0300f36f
f8d06343
f36f10a0
f8c0310c
f8d010a0
f36f20a0
f8c022cb
f8d020a0
f36f30a0
f8c033cf
f8d030a0
f36f20a0
f8c0328e
e7b920a0
68032a01
f443d10b
60023280
f4436803
60016100
20a0f8d0
7200f442
f36fe7ed
60034310
f36f6801
600121cb
20a0f8d0
2249f36f
2a01e7e1
d1136803
3100f443
68026001
5380f442
6b816003
0201f041
6b836382
0110f043
f8d06381
f44220a0
e7ca6280
4351f36f
68016003
310cf36f
6b826001
0200f36f
6b836382
1304f36f
f8d06383
f36f20a0
e7b6228a
68032a01
f443d111
60031300
f4416801
60025200
30a0f8d0
0140f043
10a0f8c0
20a0f8d0
0280f042
f36fe7a1
60035355
f36f6801
6001314d
20a0f8d0
1286f36f
20a0f8c0
20a0f8d0
12c7f36f
f8d0e78f
f44220a0
e78a3200
f0436ac3
62c10101
2a01e742
6803d116
7180f443
68026001
0380f042
69816003
3280f441
f8d06182
f04330a0
f8c00104
f8d010a0
f04220a0
e76c0208
10a0f8d0
0182f36f
10a0f8c0
20a0f8d0
02c3f36f
20a0f8c0
f36f6803
60032308
f36f6801
600111c7
f36f6982
61824210
2a01e710
6802d119
0340f042
69c16003
2280f441
69c361c2
0101f043
f8d061c1
f04220a0
f8c00302
69c130a0
3200f441
69c361c2
4180f443
f8d0e018
f36f20a0
f8c00241
69c320a0
4351f36f
69c161c3
318ef36f
680261c1
1286f36f
69c36002
4392f36f
69c161c3
0100f36f
e6d961c1
d1122a01
f4416801
60027200
f4436803
60016180
20a0f8d0
0320f042
30a0f8c0
10a0f8d0
0210f041
f8d0e707
f36f30a0
f8c01304
f8d030a0
f36f10a0
f8c01145
680210a0
2249f36f
68036002
238af36f
6d03e6af
0101f043
e6ab6501
47702001
f0002800
290b80cd
80caf200
f001e8df
3b201306
77725f4a
c2937cae
f36f6982
61820200
f36f6803
60031345
10a0f8d0
0301f041
6801e033
318ef36f
68026001
5214f36f
68036002
2100f443
e0a56001
f36f6b41
63410100
20a0f8d0
320cf36f
20a0f8c0
30a0f8d0
23cbf36f
30a0f8c0
10a0f8d0
4200f441
20a0f8c0
30a0f8d0
4380f443
6801e00b
4110f36f
68026001
22cbf36f
f8d06002
f44330a0
f8c07300
e07b30a0
f36f6802
60024251
f36f6803
6003330c
f36f6b81
63810100
f36f6b82
63821204
30a0f8d0
6380f443
6803e7e7
5355f36f
68016003
314df36f
f8d06001
f04220a0
f8c00340
f8d030a0
f04110a0
e7d40380
30a0f8d0
4351f36f
6ac2e7cf
0200f36f
e04962c2
f36f6803
60032308
f36f6801
600111c7
f36f6982
61824210
30a0f8d0
0104f043
10a0f8c0
20a0f8d0
0308f042
6803e7b3
1386f36f
69c16003
4192f36f
69c261c1
0200f36f
f8d061c2
f04330a0
f8c00102
69c210a0
3300f442
69c161c3
4280f441
e01761c2
f36f6801
60012149
f36f6802
6002228a
30a0f8d0
0120f043
10a0f8c0
20a0f8d0
0310f042
30a0f8c0
f36f6d01
65010100
47702000
47702001
460eb570
46044615
2a08b908
4620d960
f7ff2102
2d08ff23
e8dfd85a
0e05f005
2e261e16
00413936
21012000
f7ff4602
6b61f857
0144f36f
2101e03f
22002005
f84ef7ff
23016b61
2101e035
22002006
f846f7ff
23026b61
2101e02d
22002004
f83ef7ff
23036b61
2101e025
22002003
f836f7ff
23046b61
2101e01d
22002002
f82ef7ff
23056b61
6b61e015
e0122306
46012001
f7ff2200
6b61f823
e00a2307
438cf04f
06d26d9a
6a98d514
208af36f
6b616298
f3632308
63610144
06136aa2
4620d5fc
46322102
fd35f7ff
bd702000
bd702001
7001f241
b5f8bd70
4616460f
4604461d
2b06b908
4620d953
f7ff2105
6b23feb5
f443b116
e0015300
334df366
2d066323
e8dfd845
0d04f005
2d251d15
20000035
46022101
ffe2f7fe
f36f6b20
e02b0044
20052200
f7fe2101
6b20ffd9
e0212201
20062200
f7fe2101
6b20ffd1
e0192202
20042200
f7fe2101
6b20ffc9
e0112203
20032200
f7fe2101
6b20ffc1
e0092204
20022200
f7fe2101
6b20ffb9
e0012205
22066b20
0044f362
6aa16320
d5fc05c9
21054620
f7ff463a
2000fcd4
2001bdf8
e92dbdf8
460f41f0
461d4690
6018f8bd
b9184604
d8012e07
d95c2b07
21084620
fe52f7ff
f3686a23
62230300
d8522d07
f005e8df
1d150d04
38352d25
21012000
f7fe4602
6a20ff83
0044f36f
2200e033
21012005
ff7af7fe
22016a20
2200e029
21012006
ff72f7fe
22026a20
2200e021
21012004
ff6af7fe
22036a20
2200e019
21012003
ff62f7fe
22046a20
2200e011
21012002
ff5af7fe
22056a20
6a20e009
e0062206
22002001
f7fe4601
6a20ff4f
f3622207
62200044
07c86aa1
6a23d5fc
1347f366
46206223
463a2108
fc69f7ff
e8bd2000
200181f0
81f0e8bd
460fb5f8
461e4615
b9184604
d8012bff
d9652a08
210a4620
fde8f7ff
d85f2d08
f005e8df
1e160e05
39362e26
20000041
46022101
ff1cf7fe
f36f69e0
e03f0044
20052200
f7fe2101
69e0ff13
e0352201
20062200
f7fe2101
69e0ff0b
e02d2202
20042200
f7fe2101
69e0ff03
e0252203
20032200
f7fe2101
69e0fefb
e01d2204
20022200
f7fe2101
69e0fef3
e0152205
220669e0
2001e012
46012200
fee8f7fe
220769e0
f04fe00a
6d83408c
d51906da
f36f6a81
6281218a
220869e0
0044f362
6aa361e0
d5fc079b
b2f669e1
114cf366
462061e1
463a210a
fbf5f7ff
bdf82000
bdf82001
7001f241
b5f8bdf8
4615460f
4604461e
2b7fb918
2a06d801
4620d94f
f7ff2109
2d06fd73
e8dfd849
0d04f005
2d251d15
20000035
46022101
fea8f7fe
f36f69a3
e02b731f
20052200
f7fe2101
69a3fe9f
e0212201
20062200
f7fe2101
69a3fe97
e0192202
20042200
f7fe2101
69a3fe8f
e0112203
20032200
f7fe2101
69a3fe87
e0092204
20022200
f7fe2101
69a3fe7f
e0012205
220669a3
731ff362
6aa061a3
d5fc0681
f36669a1
61a14157
21094620
f7ff463a
2000fb96
2001bdf8
b538bdf8
46044615
b918461a
d8012dff
d9502907
f36f6963
61630300
d84a2907
f001e8df
1a130c04
322f2821
46012000
fe4ef7fe
f36f6960
e02d0044
21002005
fe46f7fe
22016960
2006e024
f7fe2100
6960fe3f
e01d2202
21002004
fe38f7fe
22036960
2003e016
f7fe2100
6960fe31
e00f2204
21002002
fe2af7fe
22056960
6960e008
e0052206
21002001
fe20f7fe
22076960
0044f362
6aa16160
d5fc0708
b2ed6963
134cf365
69606163
0201f040
20006162
2001bd38
e92dbd38
468841f0
461e4615
7018f8bd
28004604
2fffd060
2a08d85e
2b08d85c
2104d85a
fcb6f7ff
d00e2d01
2d02d304
2004d152
e00a2101
21012005
f7fe2200
6ba3fdeb
0343f36f
2006e007
22004629
fde2f7fe
f3656ba3
63a30343
d83b2e04
f006e8df
170f0703
6ba0001f
1048f36f
2000e01b
21014602
fdcef7fe
22016ba0
2200e011
21012003
fdc6f7fe
22026ba0
2200e009
21012002
fdbef7fe
22036ba0
6ba0e001
f3622204
63a01048
05496aa1
6aa3d5fc
d5fc051a
06436aa0
6ba2d5fc
f367b2ff
63a22250
21044620
f7ff4642
2000face
81f0e8bd
e8bd2001
b57081f0
461d460e
b9204604
d8062bff
d8042a06
6ac3e050
0300f36f
2a0662c3
e8dfd84a
0d04f002
2d251d15
20000035
46022101
fd82f7fe
f36f6ae0
e02b0044
20052200
f7fe2101
6ae0fd79
e0212201
20062200
f7fe2101
6ae0fd71
e0192202
20042200
f7fe2101
6ae0fd69
e0112203
20032200
f7fe2101
6ae0fd61
e0092204
20022200
f7fe2101
6ae0fd59
e0012205
22066ae0
0044f362
6aa162e0
d5fc0588
b2ed6ae3
134cf365
462062e3
46322107
fa6ff7ff
bd702000
bd702001
d8142905
f001e8df
0b07030b
2204110d
23007002
2104e00a
23027001
2304e006
2304e004
23057003
2301e000
20007003
79404770
79034770
71014319
79034770
0101ea23
47707101
477078c0
477070c1
47707880
f0437843
70410104
78434770
0102f043
47707041
70432306
7ec04770
7e404770
7e804770
7e004770
b5134770
46042300
f88d6800
f88d3001
f88d3002
78c13003
1001f88d
2001f89d
0308f002
b940b2d8
0001f89d
0102f000
2b00b2cb
8097f040
69a1e0f0
d0f32900
795a6823
d0ef2a00
91012100
69a168d8
9b019001
f0139801
bf180280
740a2201
69a39901
0240f010
000ff001
2201bf18
725a7218
7c1a69a3
2a01b112
e02ed16a
9a019801
2107f3c0
5042f3c2
02c1ea40
60da7a59
d15d2900
0e029801
6823701a
68d969a0
9a019101
70429901
9a0169a3
70980a08
0c1169a3
9b0170d9
0e1a69a0
68217102
68c869a3
9a019001
715a9801
9a0169a1
718b0a03
0c1269a1
9801e039
9a019901
4107f3c1
f3c00349
ea412007
0e125040
1042ea40
60d86821
920168ca
f3c19901
431002c4
7a5860d8
9901bb10
0a0a9801
69a3701a
0c019a01
69a37059
70980e10
69a06821
930168cb
9b019a01
69a170c2
0a189a01
69a17108
714b0c13
69a09901
71820e0a
69a16823
900168d8
71ca9a01
b11368a3
21014620
68214798
70c82008
6820e76c
70c22202
68e26821
f88d7e0b
2a003002
f89dd050
b9091002
47904620
0002f89d
d5030600
462068e3
47982106
1002f89d
0240f001
b118b2d0
462068e3
47982107
1002f89d
0220f001
b118b2d0
462068e3
47982108
1002f89d
0210f001
b118b2d0
462068e3
47982105
1002f89d
0208f001
b118b2d0
462068e3
47982104
1002f89d
0204f001
b118b2d0
462068e3
47982103
1002f89d
0202f001
b118b2d0
462068e3
47982102
1002f89d
d50307c9
462068e2
47902101
0001f89d
0320f000
b1c9b2d9
22206820
682370c2
69237899
1003f88d
f89db183
07c20003
4620d502
47982102
2003f89d
0102f002
b11bb2cb
46206922
47902103
0001f89d
0110f000
b13bb2cb
22106820
692370c2
4620b113
47982101
1001f89d
0040f001
b13ab2c2
21406823
692270d9
4620b112
47902104
0001f89d
d51107c3
21016823
682270d9
789068a3
0003f88d
f89db143
f0011003
b2d00240
4620b110
47982102
3001f89d
0104f003
b13ab2ca
23046820
68a270c3
4620b112
47902100
7880bd1c
0120f000
f241b2ca
2a000303
4618bf0c
47702000
4605b573
96002600
9601460c
29006169
80c1f000
f7ff6800
9001ffe8
f2419801
42980303
80bbf000
b1187c20
f0402801
e03a80a4
68e07a22
f3627a63
f3600603
08c15657
260ff361
1686f363
f0402b00
98008094
78617822
661ff362
0200ea41
98009200
ea4078a1
92002201
78e19800
4201ea40
98009200
ea407921
68286201
60869200
682a9900
93006091
79609b00
0203ea40
99009200
79e279a3
2003ea41
99009000
4302ea41
9900e063
f0417a63
92000280
2b01b12b
9800d107
0240f040
9900e002
0240f021
9b009200
ea407a20
68e30103
98009100
f4020b5a
4301417f
98009100
3247f3c3
4102ea40
98009100
095b6829
6203ea40
98009200
23006088
930068e1
00c89a00
7a60b2c3
93004313
d1322800
78219a00
2301ea42
9a009300
ea427861
93004301
78a19a00
6301ea42
99009300
6091682a
9b009000
ea4278e2
91000103
79229b00
2102ea43
9b009100
ea437962
91004102
79a29b00
6102ea43
9a009100
609a682b
98009000
ea4179e1
93000300
682b9800
7d206098
2801b128
6829d10c
704a2206
682be008
f0417859
705a0204
f241e003
e0000001
b2002000
201cbd7c
b0824770
f88d2300
f88d3006
28003007
8093f000
f0002900
7e028090
2006f88d
2006f89d
680bb91a
1307f362
f89d600b
06122006
680bd504
f3622206
600b1307
3006f89d
0240f003
b123b2d3
2207680b
1307f362
f89d600b
f0033006
b2d30220
680bb123
f3622208
600b1307
3006f89d
0210f003
b123b2d3
2205680b
1307f362
f89d600b
f0033006
b2d30208
680bb123
f3622204
600b1307
3006f89d
0204f003
b123b2d3
2203680b
1307f362
f89d600b
f0033006
b2d30202
680bb123
f3622202
600b1307
3006f89d
d50407db
2201680b
1307f362
7e42600b
f362680b
600b4317
f3627e82
600b230f
f88d7882
f89d2007
07d22007
2202d503
0303f362
7e83600b
7e82b113
d50d0612
b1137e43
06137e42
7e83d508
d9012b80
e0037e83
2a807e42
7e43d905
23016808
0003f363
6808e002
0003f36f
20006008
f241e001
b0020001
b1404770
6803b139
791a6181
0008f042
20007118
f2414770
47700001
2902b168
b152d80b
d0032901
d0032902
e0026102
e0006082
200060c2
f2414770
47700001
70032304
32fff04f
23012105
61027001
70036142
47702000
2800b510
80aff000
f0002a00
2b0080ac
80a9f000
70012104
70012105
b1197c11
f0402901
e048809c
690168d4
04c7f3c4
0107f364
68d46101
b2cc0161
f3646901
6101210f
694168dc
04c7f3c4
0107f364
68dc6141
b2cc0161
f3646941
6141210f
7a516904
2407f3c4
f004b911
e00104ef
0410f044
f3646901
6101210f
7a596944
2407f3c4
f004b911
e00104ef
0410f044
f3646941
6141210f
69017814
4117f364
69416101
f364781c
61414117
69027851
621ff361
78596102
68d4e04d
f3c46901
f3645447
61010107
690168d4
3447f3c4
210ff364
68d46101
f3c46901
f3641447
61014117
00e168d4
6901b2cc
611ff364
69016101
0e097a52
f041b112
e0010104
01fbf001
f3616902
6102621f
694268d9
5147f3c1
0207f361
68d96142
f3c16942
f3613147
6142220f
694268d9
1147f3c1
4217f361
68d96142
b2d100ca
f3616942
6142621f
7a5b6941
b1130e0a
0104f042
f002e001
694301fb
631ff361
21016143
20007001
f241bd10
bd100001
460db570
2100221c
f0074604
6868fbeb
602068ab
28006063
6828d059
1e517802
d853290f
1e5a7843
d84f2a07
1e4b7881
d84b2b03
1e428880
293fb291
f04fd846
6973468c
d4080159
6180f04f
f7fd4630
4630fa95
f7fd210c
6820fa85
70032304
68226829
79917908
f3603801
71910105
68226828
1e487881
f3607991
71911187
68226828
1e487801
f36079d1
71d10103
68226828
1e487841
f36079d1
71d11106
68286822
798079d1
11c7f360
682271d1
f0407910
71110177
49056822
20007013
f8c17010
46203188
bd70608b
bd702000
e000e100
781a6803
0104f042
68037019
f36f799a
719a0205
798b6801
1387f36f
6801718b
f36f79ca
71ca0203
79d96803
1106f36f
4b0771d9
22042100
2188f8c3
2088f8c3
60c16101
f04f6081
210c408c
ba26f7fd
e000e100
60032301
68804770
684b4770
477060c3
221f7a0b
011ff003
61016142
47702000
61c32301
220268c9
61c26181
6a0b4770
d8052b01
62022204
61c2b103
47702000
3001f241
7e0b4770
030ff003
f04f061b
62c2427f
7e096283
0713090a
20006283
7c0a4770
f0024603
28020007
6899d102
d5fc0789
07d2689a
2101d5fc
60196b98
6bcb4770
47706383
7380f44f
47706283
47706b40
7c0cb510
0407f004
dc182c02
f04f2c01
f04f0320
d0040240
d00a2c02
62c262c3
6283e00b
62c2231f
7c0a62c3
628108d1
6282e003
694962c3
20006301
f241bd10
bd103001
2a016a4a
2380d80c
6283b10a
62c3e000
f0126b42
d1fb0304
624169c9
47704618
3001f241
7b034770
0101f043
47707301
f0237b03
73010101
69c34770
0107f001
0203ea41
477061c2
b2c06940
68034770
60014319
79034770
0108f043
47707101
f0437903
71010102
79034770
0101f043
47707101
f0437a03
72010108
7a034770
0102f043
47707201
f0437a03
72010101
00004770
460db5f8
46044617
2931b1f8
2601d820
f3f3fbb6
707af44f
f0064358
4601ff93
f007480d
f007f89b
b2c0f9d1
f4410101
f10562a0
4332458c
f5052000
61e24560
626060e6
703b782b
f640bdf8
bdf82003
2001f640
bf00bdf8
42280000
460eb5f8
46044617
2931b1f8
2501d820
f3f3fbb5
707af44f
f0064358
4601ff65
f007480d
f007f86d
b2c0f9a3
f4410101
f10662a0
432a468c
4660f506
60e561e2
88336265
803b2000
f640bdf8
bdf82003
2001f640
bf00bdf8
42280000
b1e0b510
d81d2931
d81e2a07
60c42406
1142ea41
2204240b
7300f443
60016084
63436042
054b6981
220ad5fc
60422301
68c16043
0202f001
200060c2
f640bd10
bd102003
2001f640
f640bd10
bd102002
2931b198
69c3d814
0301f043
f44161c3
23014100
60c36101
04096941
2300d5fc
694060c3
46187010
f6404770
47702003
2001f640
00004770
b087b530
f89d2b01
d8134028
93032300
9b030080
d25e428b
9b039c03
f103009b
f5035310
581b23c0
3024f842
33019b03
e7ee9303
d1122b02
93032300
9b030080
d248428b
9c039b03
f10400a4
f5045410
582424c0
9b0354d4
93033301
2b03e7ef
0080d139
2300b32c
9b049304
d232428b
006c9d04
9b059405
f105005d
f5045410
5a1d23c0
f88db2ec
9b054008
005d4c13
5a1d192b
f88db2ec
9b044004
5004f89d
4008f89d
2405ea44
4013f822
33019b04
9403e7da
428b9b03
9b03d20d
00a49c03
5410f104
24c0f504
f8225824
9b034013
93033301
b007e7ee
bf00bd30
24060002
b085b530
93032300
9b030092
d226428b
f3448804
b2ab2507
3004f8ad
4b02f830
f88db2a5
f89d5003
b25c3003
4008f8ad
006b9d03
005cb29b
5510f104
24c0f505
5008f8bd
52a5b2ad
4b06005c
f8bd18e3
b2a44004
9b03529c
93033301
b005e7d5
bf00bd30
24060002
1181ea40
ea414b02
61da4202
bf004770
24070000
4b0db530
f0046a1c
2a03647c
e8dfd812
020af002
f4440805
e0047480
7400f444
f444e001
f0447440
ea440401
ea404000
62192181
bf00bd30
24070000
41f0e92d
b2d1460e
46154c16
460a4607
46982000
ffccf7ff
61a3231f
46294638
f7ff2200
4630ff91
f44f4629
f7ff7200
6861ff8b
010cf36f
68a06061
7200f44f
000cf362
68e160a0
6380f44f
010cf363
60e1208f
20006020
46424601
41f0e8bd
bfb0f7ff
24070000
41f0e92d
b2d1460e
46154c16
460a4607
46982000
ff98f7ff
61a3231f
46294638
f7ff2200
4630ff5d
f44f4629
f7ff7200
6861ff57
010cf36f
68a06061
7200f44f
000cf362
68e160a0
6380f44f
010cf363
60e12093
20006020
46424601
41f0e8bd
bf7cf7ff
24070000
460eb5f8
4c16b2d1
46074615
2000460a
ff66f7ff
61a32319
46294638
f7ff2200
4630ff2b
f44f4629
f7ff7200
6860ff25
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002195
220160e3
46016021
40f8e8bd
bf4af7ff
24070000
460eb5f8
4c16b2d1
46074615
2000460a
ff34f7ff
61a32319
46294638
f7ff2200
4630fef9
f44f4629
f7ff7200
6860fef3
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002195
220260e3
46016021
40f8e8bd
bf18f7ff
24070000
460eb5f8
4c16b2d1
46074615
2000460a
ff02f7ff
61a32319
46294638
f7ff2200
4630fec7
f44f4629
f7ff7200
6860fec1
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002195
220360e3
46016021
40f8e8bd
bee6f7ff
24070000
b570b2d1
46064c10
20004615
f7ff460a
2319fed1
463061a3
22004629
fe96f7ff
f36f6860
6060000c
f44f68e1
f3627200
2000010c
f24060e1
46011357
60232203
4070e8bd
bec0f7ff
24070000
60828001
47706043
60828001
47706043
60828001
47706043
60828001
47706043
60828001
4a036819
611160c3
6153685b
bf004770
24070000
60828001
4a036819
611160c3
6153685b
bf004770
24070000
60828001
1000f9b3
60c34a03
f9b36111
61533002
bf004770
24070000
fb92b510
fb01f4f1
b9322214
9b026043
80447001
46106083
20fee000
bd10b240
f4436803
60016180
b5104770
f1010089
f5035310
230021c0
d0054293
4023f850
f8413301
e7f74b04
b510bd10
d8252b03
f003e8df
02091010
f1010089
f5035310
230021c0
008ce012
5110f104
21c0f501
e0032300
4010e8bd
bfd7f7ff
d0044293
330156c4
4b04f841
bd10e7f8
d0054293
4013f930
f8413301
e7f74b04
0000bd10
460eb5f8
4c17b2d9
460a4607
461d2000
fe24f7ff
61a3231f
21004638
2302462a
ffc3f7ff
462a4630
f44f2302
f7ff7100
6860ffbc
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
2000218f
460260e3
46016021
40f8e8bd
be06f7ff
24070000
460eb5f8
4c17b2d9
460a4607
461d2000
fdf0f7ff
61a3231f
21004638
2303462a
ff8ff7ff
462a4630
f44f2303
f7ff7100
6860ff88
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
2000218f
460260e3
46016021
40f8e8bd
bdd2f7ff
24070000
460eb5f8
4c17b2d9
460a4607
461d2000
fdbcf7ff
61a3231f
21004638
2302462a
ff5bf7ff
462a4630
f44f2302
f7ff7100
6860ff54
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002193
460260e3
46016021
40f8e8bd
bd9ef7ff
24070000
460eb5f8
4c17b2d9
460a4607
461d2000
fd88f7ff
61a3231f
21004638
2303462a
ff27f7ff
462a4630
f44f2303
f7ff7100
6860ff20
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002193
460260e3
46016021
40f8e8bd
bd6af7ff
24070000
460eb5f8
4c17b2d9
460a4607
461d2000
fd54f7ff
61a32319
21004638
2302462a
fef3f7ff
462a4630
f44f2302
f7ff7100
6860feec
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002195
460260e3
46016021
40f8e8bd
bd36f7ff
24070000
460eb5f8
4c17b2d9
460a4607
461d2000
fd20f7ff
61a32311
21004638
2303462a
febff7ff
462a4630
f44f2303
f7ff7100
6860feb8
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002195
460260e3
46016021
40f8e8bd
bd02f7ff
24070000
460db570
4c11b2c9
460a4606
f7ff2000
2319fced
463061a3
462a2100
f7ff2302
6860fe8c
000cf36f
68e16060
7200f44f
010cf362
60e12000
1357f240
46024601
e8bd6023
f7ff4070
bf00bcdb
24070000
460db570
4c11b2c9
460a4606
f7ff2000
2311fcc5
463061a3
462a2100
f7ff2303
6860fe64
000cf36f
68e16060
7200f44f
010cf362
60e12000
1357f240
46024601
e8bd6023
f7ff4070
bf00bcb3
24070000
41f0e92d
460f9e06
4690b2f1
460a4604
461d7800
fc9af7ff
46384b1a
8018f8c3
4631b155
f7ff2200
68a0fc5d
f44f8821
f7ff7200
e00bfc57
46324629
f7ff2303
68a0fe2c
f44f8822
23037100
fe25f7ff
6841480c
010cf36f
68836041
7200f44f
030cf362
68c16083
6380f44f
010cf363
60c12203
20006002
462a4601
41f0e8bd
bc6ef7ff
24070000
41f0e92d
46884c18
4605b2d9
4617461e
460a7800
fc56f7ff
21004640
23024632
f7ff61a7
68a8fdf6
2302882a
7100f44f
fdeff7ff
f36f6863
6063030c
f44f68a0
f3627200
60a0000c
f44f68e1
f3636380
2003010c
602060e1
46012000
e8bd4602
f7ff41f0
bf00bc39
24070000
41f0e92d
b2d9460f
46044690
7800460a
5018f89d
f7ff461e
4b1bfc1f
f8c34638
b1558018
22004631
fbe2f7ff
882168a0
7200f44f
fbdcf7ff
4629e00b
23034632
fdb1f7ff
882268a0
7100f44f
f7ff2303
480dfdaa
f36f6842
6042020c
f44f6883
f3617100
6083030c
f44f68c2
f3636380
2105020c
600160c2
46012000
e8bd462a
f7ff41f0
bf00bbf3
24070000
43f8e92d
78044699
f89d8843
435c6020
b2e04605
46174688
4602b2d1
fbd6f7ff
b1564640
22004639
fb9cf7ff
46216868
7200f44f
fb96f7ff
4631e00b
2303463a
fd6bf7ff
f44f6868
46227100
f7ff2303
4c10fd64
9018f8c4
f36f6860
6060000c
f44f68a1
f3627200
60a1010c
f44f68e3
f3606080
21c7030c
602160e3
6a23782a
5082ea43
20006220
46324601
43f8e8bd
bba6f7ff
24070000
460db5f8
882a884f
88068841
d12f428a
b2d34c19
61e32111
437261a1
68402303
7100f44f
fd2df7ff
886a882b
435a6868
6180f44f
f7ff2303
6860fd24
7200f44f
000cf362
68a16060
6380f44f
010cf363
68e060a1
62c0f44f
000cf362
60e02199
60212200
46394630
fb6ef7ff
bdf82000
0001f242
bf00bdf8
24070000
460eb5f8
4c16b2d1
46074615
2000460a
fb52f7ff
61a3231f
21004638
f7ff462a
4630fce2
f44f462a
f7ff7100
6860fcdc
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
2000218f
460260e3
46016021
40f8e8bd
bb36f7ff
24070000
460eb5f8
4c16b2d9
460a4607
461d2000
fb20f7ff
61a3231f
21004638
f7ff462a
4630fcb0
f44f462a
f7ff7100
6860fcaa
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
2000218f
460260e3
46016021
40f8e8bd
bb04f7ff
24070000
41f0e92d
b2d1460e
46154c16
460a4607
46982000
faecf7ff
61a3231f
21004638
f7ff462a
4630fc7c
f44f462a
f7ff7100
6861fc76
010cf36f
68a06061
7200f44f
000cf362
68e160a0
6380f44f
010cf363
60e1208f
20006020
46424601
41f0e8bd
bad0f7ff
24070000
41f0e92d
b2d1460e
46154c16
460a4607
46982000
fab8f7ff
61a3231f
21004638
f7ff462a
4630fc48
f44f462a
f7ff7100
6861fc42
010cf36f
68a06061
7200f44f
000cf362
68e160a0
6380f44f
010cf363
60e1208f
20006020
46424601
41f0e8bd
ba9cf7ff
24070000
460eb5f8
4c16b2d1
46074615
2000460a
fa86f7ff
61a3231f
21004638
f7ff462a
4630fc16
f44f462a
f7ff7100
6860fc10
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002193
460260e3
46016021
40f8e8bd
ba6af7ff
24070000
43f8e92d
f89d4c18
46889020
461eb2d9
46174605
460a7800
fa50f7ff
21004640
61a74632
fbe1f7ff
882a68a8
7100f44f
fbdbf7ff
f36f6863
6063030c
f44f68a0
f3627200
60a0000c
f44f68e1
f3636380
2005010c
602060e1
46012000
e8bd464a
f7ff43f8
bf00ba35
24070000
43f8e92d
f89d4c18
46889020
461eb2d9
46174605
460a7800
fa1af7ff
21004640
61a74632
fbabf7ff
882a68a8
7100f44f
fba5f7ff
f36f6863
6063030c
f44f68a0
f3627200
60a0000c
f44f68e1
f3636380
2005010c
602060e1
46012000
e8bd464a
f7ff43f8
bf00b9ff
24070000
41f0e92d
4604461d
78008843
f89d9e06
4358801c
460fb2c0
b2e94602
f9e2f7ff
21004638
f7ff462a
4b10fb74
6859619e
010cf36f
68986059
7200f44f
000cf362
68d96098
6080f44f
010cf360
6a1a60d9
ea427821
62185081
200022c7
4601601a
e8bd4642
f7ff41f0
bf00b9c7
24070000
fb92b538
fb01f5f1
b92c2415
9b046043
80457001
e0006083
684024fe
7100f44f
fb3ff7ff
bd38b260
fb92b538
fb01f5f1
b92c2415
9b046043
80457001
e0006083
684024fe
7100f44f
fb2bf7ff
bd38b260
41f0e92d
4604461d
78008843
f89d9e06
4358801c
460fb2c0
b2e94602
f982f7ff
21004638
f7ff462a
4b10fb14
6859619e
010cf36f
68986059
7200f44f
000cf362
68d96098
6080f44f
010cf360
60d922c7
6a18601a
ea407821
20005281
4601621a
e8bd4642
f7ff41f0
bf00b967
24070000
460eb5f8
4c16b2d9
460a4607
461d2000
f950f7ff
61a3231f
21004638
f7ff462a
4630fae0
f44f462a
f7ff7100
6860fada
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002193
460260e3
46016021
40f8e8bd
b934f7ff
24070000
41f0e92d
b2d1460e
46154c16
460a4607
46982000
f91cf7ff
61a3231f
21004638
f7ff462a
4630faac
f44f462a
f7ff7100
6861faa6
010cf36f
68a06061
7200f44f
000cf362
68e160a0
6380f44f
010cf363
60e12093
20006020
46424601
41f0e8bd
b900f7ff
24070000
41f0e92d
b2d1460e
46154c16
460a4607
46982000
f8e8f7ff
61a3231f
21004638
f7ff462a
4630fa78
f44f462a
f7ff7100
6861fa72
010cf36f
68a06061
7200f44f
000cf362
68e160a0
6380f44f
010cf363
60e12093
20006020
46424601
41f0e8bd
b8ccf7ff
24070000
41f0e92d
460f4c17
461db2d9
46164680
460a2000
f8b4f7ff
21004640
61a6462a
fa45f7ff
462a4638
7100f44f
fa3ff7ff
f36f6863
6063030c
f44f68a0
f3627200
60a0000c
f44f68e1
f3636380
2095010c
602060e1
46012000
e8bd4602
f7ff41f0
bf00b899
24070000
460eb5f8
4c16b2d9
460a4607
461d2000
f882f7ff
61a32301
21004638
f7ff462a
4630fa12
f44f462a
f7ff7100
6860fa0c
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002195
460260e3
46016021
40f8e8bd
b866f7ff
24070000
41f0e92d
460f4c17
4615b2d1
460a4680
26012000
f84ef7ff
21004640
61a6462a
f9dff7ff
462a4638
7100f44f
f9d9f7ff
f36f6863
6063030c
f44f68a0
f3627200
60a0000c
f44f68e1
f3636380
2095010c
602060e1
46012000
e8bd4632
f7ff41f0
bf00b833
24070000
41f0e92d
460f4c17
461db2d9
46164680
460a2000
f81af7ff
21004640
61a6462a
f9abf7ff
462a4638
7100f44f
f9a5f7ff
f36f6863
6063030c
f44f68a0
f3627200
60a0000c
f44f68e1
f3636380
2095010c
602060e1
46012000
e8bd2201
f7fe41f0
bf00bfff
24070000
41f0e92d
460f4c17
461db2d9
46164680
460a2000
ffe6f7fe
21004640
61a6462a
f977f7ff
462a4638
7100f44f
f971f7ff
f36f6863
6063030c
f44f68a0
f3627200
60a0000c
f44f68e1
f3636380
2095010c
602060e1
46012000
e8bd2202
f7fe41f0
bf00bfcb
24070000
460eb5f8
4c16b2d9
460a4607
461d2000
ffb4f7fe
61a32301
21004638
f7ff462a
4630f944
f44f462a
f7ff7100
6860f93e
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002195
220260e3
46016021
40f8e8bd
bf98f7fe
24070000
41f0e92d
460f4c17
461db2d9
46164680
460a2000
ff80f7fe
21004640
61a6462a
f911f7ff
462a4638
7100f44f
f90bf7ff
f36f6863
6063030c
f44f68a0
f3627200
60a0000c
f44f68e1
f3636380
2095010c
602060e1
46012000
e8bd2203
f7fe41f0
bf00bf65
24070000
460eb5f8
4c16b2d9
460a4607
461d2000
ff4ef7fe
61a32311
21004638
f7ff462a
4630f8de
f44f462a
f7ff7100
6860f8d8
000cf36f
68a16060
7200f44f
010cf362
68e360a1
6080f44f
030cf360
20002195
220360e3
46016021
40f8e8bd
bf32f7fe
24070000
b570b2d1
46064c10
20004615
f7fe460a
2301ff1d
463061a3
462a2100
f8adf7ff
f36f6860
6060000c
f44f68e1
f3627200
2000010c
f24060e1
46011357
60232203
4070e8bd
bf0cf7fe
24070000
460db570
4c10b2c9
460a4606
f7fe2000
2301fef7
463061a3
462a2100
f887f7ff
f36f6860
6060000c
f44f68e1
f3627200
2000010c
f24060e1
46011357
60234602
4070e8bd
bee6f7fe
24070000
460db570
4c10b2c9
460a4606
f7fe2000
2309fed1
463061a3
462a2100
f861f7ff
f36f6860
6060000c
f44f68e1
f3627200
2000010c
f24060e1
46011357
60234602
4070e8bd
bec0f7fe
24070000
460db5f8
882b884f
88068841
d12d428b
b2d94c18
61a261e1
fb036840
f44ff206
f7ff7100
882bf838
6868886a
f44f435a
f7ff6180
6860f830
7200f44f
000cf362
68a16060
6380f44f
010cf363
68e060a1
62c0f44f
000cf362
60e02199
60212200
46394630
fe8af7fe
bdf82000
0001f242
bf00bdf8
24070000
460db5f8
882a884f
88068841
d12d428a
b2d34c18
61e32101
437261a1
f44f6840
f7fe7100
882bfffc
6868886a
f44f435a
f7fe6180
6860fff4
7200f44f
000cf362
68a16060
6380f44f
010cf363
68e060a1
62c0f44f
000cf362
60e02199
60212200
46394630
fe4ef7fe
bdf82000
0001f242
bf00bdf8
24070000
43f8e92d
4c179e08
b2f14688
46174605
460a7800
f7fe4699
4640fe2f
46322100
f7fe61a7
68a8ffc0
f44f882a
f7fe7100
6861ffba
010cf36f
68a06061
7300f44f
000cf363
68e260a0
6180f44f
020cf361
60e22003
20006020
464a4601
43f8e8bd
be14f7fe
24070000
43f8e92d
4c179e08
b2f14688
46174605
460a7800
f7fe4699
4640fdfb
46322100
f7fe61a7
68a8ff8c
f44f882a
f7fe7100
6861ff86
010cf36f
68a06061
7300f44f
000cf363
68e260a0
6180f44f
020cf361
60e22003
20006020
464a4601
43f8e8bd
bde0f7fe
24070000
9b04b538
b2dd4c0e
61e501ad
612161a2
2100461a
f7fe2303
6860ff6e
000cf36f
68e16060
7200f44f
010cf362
60e12000
4601238d
60234602
4038e8bd
bdbef7fe
24070000
9b04b538
b2dd4c0e
61e501ad
612161a2
2100461a
ff3df7fe
f36f6860
6060000c
f44f68e1
f3627200
2000010c
238d60e1
46024601
e8bd6023
f7fe4038
bf00bd9d
24070000
4c0fb538
b2d3461d
61e3019b
61a32315
21006121
ff1bf7fe
f36f6861
6061010c
f44f68e0
f3627200
60e0000c
238d2000
462a4601
e8bd6023
f7fe4038
bf00bd7b
24070000
4c1bb573
b2d3461e
4611460d
2319019a
61a361e2
f7fe2200
1228fd2d
f88db2ed
f88d0003
f89d5002
b24a1003
2004f8ad
3002f89d
f8adb258
f8bd0006
f8bd1004
b2932006
4001ea43
68616120
010cf36f
68e26061
7300f44f
020cf363
60e2208d
20006020
46324601
fd42f7fe
bf00bd7c
24070000
4c0fb538
b2d3461d
61e3019b
61a32301
21006121
febff7fe
f36f6861
6061010c
f44f68e0
f3627200
60e0000c
238d2000
462a4601
e8bd6023
f7fe4038
bf00bd1f
24070000
b2d3b510
019b4c0d
61a161e3
f7fe2100
6860fea0
000cf36f
68e16060
7200f44f
010cf362
60e12000
1357f240
22034601
e8bd6023
f7fe4010
bf00bcff
24070000
4c0eb538
01adb2dd
61a261e5
461a6121
f7fe2100
6863fe7e
030cf36f
68e06063
7200f44f
000cf362
218960e0
60212000
46014602
4038e8bd
bcdef7fe
24070000
b2dab510
01924c0e
221f61e2
612161a2
2100461a
f7fe2302
6863fe6c
030cf36f
68e06063
7100f44f
000cf361
228960e0
60222000
46024601
4010e8bd
bcbcf7fe
24070000
b2dab510
01924c0e
221f61e2
612161a2
2100461a
f7fe2303
6863fe4a
030cf36f
68e06063
7100f44f
000cf361
228960e0
60222000
46024601
4010e8bd
bc9af7fe
24070000
b2dab510
01924c0e
221f61e2
612161a2
2100461a
fe19f7fe
f36f6863
6063030c
f44f68e0
f3617100
60e0000c
20002289
46016022
e8bd4602
f7fe4010
bf00bc79
24070000
4c0fb538
b2d3461d
61e3019b
61a3231f
21006121
fdf7f7fe
f36f6861
6061010c
f44f68e0
f3627200
60e0000c
23892000
462a4601
e8bd6023
f7fe4038
bf00bc57
24070000
4c1bb573
b2d3461e
4611460d
231f019a
61a361e2
f7fe2200
1228fc09
f88db2ed
f88d0003
f89d5002
b24a1003
2004f8ad
3002f89d
f8adb258
f8bd0006
f8bd1004
b2932006
4001ea43
68616120
010cf36f
68e26061
7300f44f
020cf363
60e22089
20006020
46324601
fc1ef7fe
bf00bd7c
24070000
4c0fb538
b2d3461d
61e3019b
61a3231f
21006121
fd9bf7fe
f36f6861
6061010c
f44f68e0
f3627200
60e0000c
23892000
462a4601
e8bd6023
f7fe4038
bf00bbfb
24070000
4c0fb538
b2d3461d
61e3019b
61a3231f
21006121
fd79f7fe
f36f6861
6061010c
f44f68e0
f3627200
60e0000c
238b2000
462a4601
e8bd6023
f7fe4038
bf00bbd9
24070000
4c0fb538
460db2d3
231f0199
61a361e1
23032100
fd67f7fe
68606125
000cf36f
68e16060
7200f44f
010cf362
60e12000
4601238b
60234602
4038e8bd
bbb6f7fe
24070000
b2dab573
5018f89d
460e4c1e
221f0191
61a261e1
4619b1e5
f7fe2200
1233fb67
f88db2f6
f88d3003
f89d6002
b2410003
1004f8ad
2002f89d
f8adb253
f8bd3006
f8bd0004
b28a1006
4300ea42
e0056123
4629461a
f7fe2303
6126fd24
68414809
010cf36f
68c26041
7300f44f
020cf363
60c2218b
20006001
462a4601
fb74f7fe
bf00bd7c
24070000
4c0fb538
b2d3461d
61e3019b
61a3231f
21006121
fcf1f7fe
f36f6861
6061010c
f44f68e0
f3627200
60e0000c
238b2000
462a4601
e8bd6023
f7fe4038
bf00bb51
24070000
4c0eb538
01adb2dd
61a261e5
461a6121
f7fe2100
6863fcd0
030cf36f
68e06063
7200f44f
000cf362
218d60e0
60212000
46014602
4038e8bd
bb30f7fe
24070000
9b04b538
b2dd4c0e
61e501ad
612161a2
2100461a
f7fe2302
6860fcbe
000cf36f
68e16060
7200f44f
010cf362
60e12000
4601238d
60234602
4038e8bd
bb0ef7fe
24070000
8a1a6803
42c0f422
6803821a
f0428a1a
821a0201
8a1a6803
0103f001
42c0f422
3141ea42
68008219
f0238a03
82020201
68024770
f4236913
f02151ff
f043031f
61110101
6a026800
d5fc0553
68034770
47706a18
d803297f
20006803
47706299
1001f241
297f4770
6803d803
62592000
f2414770
47701001
6a986803
68034770
f4228b9a
83997180
8b836800
7200f423
20008382
203c4770
b5f04770
0343eb01
42942400
d029b2a6
6a2f6805
d42507f9
f0617e29
762e067f
6a876805
7e2f7879
060ff001
010ff027
76294331
f8336805
f8c56014
68066080
f4276937
6a8741ff
057ff021
f0457839
ea450502
61353541
6a2e6805
d4fc07f6
e7d23401
bdf04630
eb01b5f0
24000343
b2a64294
6805d01e
07f96a2f
8aa9d41a
7680f441
680582ae
f4216929
f02646c0
6a860103
f0417836
ea410184
61293146
6a2e6805
d4fc0636
1080f8d5
1014f823
e7dd3401
bdf04630
2400b5f0
b2a64294
6805d030
f0176a2f
d12b0f01
f0667e2e
762f077f
8aae6805
6780f426
680582af
78776a86
f0077e2e
f026070f
433e060f
762e18cf
68055d3e
6080f8c5
69356806
47fff425
057ff027
783f6a87
0502f045
3547ea45
68066135
f0156a35
d1fb0f01
e7cb3401
bdf04630
2400b5f0
b2a64294
6805d01f
f0176a2f
d11a0f01
f4268aae
82af7780
692e6805
47c0f426
0603f027
0784f046
78366a86
3646ea47
6805612e
06366a2e
f8d5d4fc
18cd6080
3401552e
4630e7dc
2300bdf0
3035f880
3036f880
b5104770
78196a83
d8112903
22016803
fa02695c
ea24f101
61590101
6a806803
78006959
f200fa02
615a430a
bd102000
1001f241
6a83bd10
2a03781a
6803d809
69592001
f202fa00
0102ea21
20006159
f2414770
47701001
6a826a43
b5106859
fbb16854
f013f3f4
d1010f01
e0046094
fbb14c06
4361f1f3
68006091
0247f3c3
1038f890
2038f880
bf00bd10
000f4240
d80a2903
f001e8df
08060402
47706082
477060c2
47706102
47706142
6804b530
f0017e25
f025010f
4329050f
68017621
2080f8c1
690a6801
42fff422
027ff022
0202f042
3343ea42
6800610b
07cb6a01
bd30d4fc
6804b510
f4236923
f02343ff
f043037f
f0210304
430b0107
3242ea43
68006122
061a6a03
f8d0d4fc
bd100080
d80b2a01
b11a6803
f0417819
e0020002
f022781a
70180002
47702000
1001f241
b5104770
07a04604
6848d173
d0712800
6261680b
60606023
f442889a
80986000
6a616823
78197c4a
0001f002
0201f021
701a4302
6a606823
7a81889a
0001f001
0101f022
80994301
68206a63
7c1a7a99
ffc6f7ff
68216a60
b1927a02
f042888a
808b0302
88816820
0204f041
68238082
f0408898
80990108
889a6823
0110f042
888be011
0002f023
68218088
f022888a
808b0304
88816820
0208f021
68238082
f0208898
80990110
68216a63
b1287a58
ea6f8a0a
ea6f4342
e0024053
04538a0a
82080c58
6a616820
8b817b8a
030ff002
020ff021
8382431a
6a636820
7b198b82
030ff001
01f0f022
1303ea41
46208383
2000bd10
0000bd10
f012690a
e92d5300
460441f0
d008460d
2b0068c3
4798d02f
20206821
e8bd6308
f01281f0
6ac66880
d0096849
d21e428e
69852201
47a84911
62e21982
81f0e8bd
d20e428e
46332201
68296987
686b47b8
42981980
d30e62e0
b14368e3
46294620
f8844798
f8848035
e8bd8036
f88481f0
f8843035
e8bd3036
bf0081f0
003008c4
f013690b
b5f75380
460d4604
6903d006
4798b30b
22026821
e01c630a
68ca6b06
429669c7
2202d309
2034f880
0106f10d
47b82201
63201980
6889e00d
46332201
68e947b8
42881980
d3046320
b1136923
46294620
bdfe4798
6803b538
6ada6a05
07d26a1a
d40e4604
784a6a81
6a03619a
685a6ac1
d3064291
f7ff7d99
6963fd7a
46206a21
f8944798
28010035
6869d107
682ab909
4620b11a
f7ff4629
6a23ff71
68d96b20
d2054288
b11a689a
46294620
ffa6f7ff
6ae06a23
42886859
2200d311
2035f884
46207d99
fd3af7ff
203f6823
46296318
462068a2
6a214790
2304f241
6a20828b
68c26b21
bf244291
2205f241
bd388282
460db538
b9104604
1001f241
2900bd38
62a1d0fa
1e59784b
d8f5290f
2a00686a
f7ffd0f2
6aa0fe4b
b11b7883
f7ff4620
e016fe1a
8a8a6821
0010f022
68238288
f0218a99
829a0220
8a836820
0140f023
68208281
f0228a82
82830380
f7ff4620
6820fe1c
68ca6aa1
05938a01
52fff421
0118f022
43d3ea41
78688203
d9032808
49054b04
e00261a3
49054a04
61e161a2
bd382000
0030a697
0030a6fd
0030a74d
0030a7bd
460db538
28004604
2900d07e
7d8bd07c
d9032b03
1001f241
bd388288
68216908
f0108a8a
bf146f00
5280f442
5280f422
2000828a
1303f241
62252101
f88482ab
f8840034
f8841035
692a0036
00936320
d52762e0
7e186823
017ff060
68237619
f4228a9a
82986080
6aa16823
7e19784a
000ff002
020ff021
761a4302
69186823
f0406919
f4210202
f02040c0
ea420105
6aa20001
ea407811
61183041
462068e3
47984629
00d0692a
6821d515
f4208a88
828b7380
69026820
41c0f422
f0216aa2
f0430301
78130104
3143ea41
69226101
46294620
69284790
da092800
f7ff4620
f9b5feef
f2411014
42911203
e009d0f6
d5070041
68236aa1
619a784a
23126820
3080f8c0
bd382000
1001f241
2028bd38
20244770
68434770
47708099
f8936843
f042206c
f8830001
4770006c
f8936843
f022206c
f8830001
4770006c
dc092907
7b1a6843
0107f001
0007f022
73194301
47702000
4001f240
68434770
61192000
68434770
b2c06918
29014770
6843d804
61190209
47702000
4001f240
1e8b4770
d8072bfd
b2c96840
2094f890
1094f880
47702000
4001f240
00004770
1e4a4b05
d803429a
67c16840
47702000
4001f240
bf004770
00fffffe
29016843
bf0c6b19
ea21430a
631a0202
68434770
7200f44f
4770611a
881a6843
0020f042
47708018
d1052901
f8d16841
f3c22080
47700040
6843b929
0080f8d3
0001f000
f2404770
47704001
6f186843
47704008
6843b510
206cf893
0001f022
006cf883
790a7808
d1042802
00a0f893
20a0f883
2803e005
f893bf04
f88300a4
881820a4
0240f040
8818801a
0220f040
7848801a
d8212807
2a07788a
78cad81e
d81b2a01
28037808
0314d818
809ab2a2
7808881c
0442f360
881a801c
0001f042
20008018
784a6318
403cf893
203cf883
f893788a
f8831038
bd102038
4001f240
b149bd10
f44f2300
61c16281
6203608a
83cb838b
47704610
4001f240
68434770
206cf893
0001f022
006cf883
f36f881a
801a0200
891a8888
0209f360
8818811a
1086f36f
784a8018
d8242a07
28077888
78cad821
d81e2a01
28037808
881ad81b
0020f042
881a8018
f36078c8
801a02c3
881a7808
0242f360
6888801a
784a6318
003cf893
203cf883
f8937888
f8831038
20000038
f2404770
47704001
460db537
0103f010
d1104604
f0042224
6868ff97
6060682b
f8906023
f022206c
f8800101
6c03106c
93014620
2000e000
b537bd3e
f010460d
46040103
2228d10a
ff7ef004
682b6868
60236060
46206c01
e0009101
bd3e2000
b5102b02
2b03d00e
2b01d015
2905d11b
6843d902
82998a9c
d9142a07
8b016840
bd108302
bf842905
83996843
d90a2a07
840a6841
2905bd10
6843bf84
2a078499
6843bf84
bd10851a
6182b909
29014770
6102d101
29024770
6142d101
29034770
6082d101
29044770
60c2bf08
b9094770
47706082
d1012901
477060c2
d1012902
47706102
d1012903
47706142
bf082904
47706182
6842b530
8d9169c4
f001b289
b2ad0540
4603b08b
d0562d00
0080f8d2
7f80f5b0
d817d042
d0392808
2802d807
2804d032
2801d032
210fd144
2820e041
d803d030
d13d2810
e03a2113
d02b2840
d1372880
e0342116
3f00f5b0
d80ad02c
5f80f5b0
f5b0d024
d0233f80
6f00f5b0
211ad128
f5b0e025
d01f2f00
f5b0d804
d11f2f80
e01c2121
1f80f5b0
f5b0d018
d1170f00
e0142124
e0122110
e0102111
e00e2112
e00c2114
e00a2115
e0082117
e006211b
e004211f
e0022120
e0002122
60a12123
92016c12
f401e11f
b2ad4580
210eb125
6c126201
e0379202
5500f401
b125b2ad
6201210d
92036c12
f401e02e
b2ad6500
210bb13d
62016852
f0026e92
92040201
f401e022
b2ad6580
210ab13d
62016852
f0026e52
92050201
f401e016
b2ad7500
2109b13d
62016852
f0026e12
92060201
f401e00a
b2ad7580
2108b175
62016852
f0026dd2
92070201
60a1689b
f0002b00
462180e3
e0df4798
0004f001
b308b280
8a617e60
b191b198
1088f892
0001f041
0088f882
0090f892
f0037ee3
f0200107
430b0307
3090f882
76622200
b121e09d
6f106861
d5fc0700
f44fe08f
61107000
e0b96219
0010f001
2800b280
8096f000
8a217e20
b319b118
76212100
b1f9e01e
68202901
d10f8c99
f4405c40
61107000
8a211c4a
1e48849a
69228220
f0402a00
621a809b
e08f68da
8a105c45
00fff020
82104328
849a1c4a
1e598a23
e08b8221
29008a61
6aa0d063
d12b2801
21027e60
62a12801
f892d10f
f0411088
f8820001
7ee10088
0007f001
1090f892
0107f021
f8824301
88101090
0120f040
f8928011
f020006c
f8820101
8aa0106c
f8928090
f041106c
f8820001
8ae1006c
7000f441
6111b281
8a617e60
2900b1a0
2901d054
f44fbf0c
f44f7140
61117180
2a076ae2
699ad104
4618b112
47904621
1c596ae3
e01862e1
d03f2900
d1072901
7140f44f
68616111
07006f10
e006d5fc
7080f44f
68616110
07006f10
6910d5fc
54888cda
1c488cd9
8a6384d8
82621e5a
6219e024
2a017e62
699abf0c
e015691a
d50707c8
21006850
6c426219
0001f002
e0099008
0102f001
b160b288
68502101
6c826219
9209400a
689a60a1
4618b132
47904621
f240e002
621a4212
bd30b00b
4605b5f8
2900460c
8097f000
6f1e6843
0601f016
4212f240
608ad002
bdf84610
61e96f1f
4707f240
6202608f
84868a0a
b34a84c6
2a017e0a
206cf893
0201f022
206cf883
809a8a8a
206cf893
0201f042
206cf883
611a8aca
f893d111
f0466088
f8830202
f8932088
7e8e208c
0207f022
0607f006
f8834332
6943208c
f8d3e02d
07c00080
e044d4fb
b3728a4a
2a017e4a
206cf893
0201f022
206cf883
809a8a8a
206cf893
0201f042
206cf883
f4428aca
b2927280
d113611a
6088f893
0201f046
2088f883
2090f893
f0227ece
f0060207
43320607
2090f883
b1d36983
e0184798
1080f8d3
d4fb07c9
f893e013
f020006c
f8830101
8aa2106c
f893809a
f040006c
f8830101
8ae2106c
f8d3611a
07c20080
686bd4fb
6b1969e0
0200ea41
68e3631a
d40107db
bdf868a0
f24068a1
42814007
4628d1f8
fdd6f7ff
f240e7f6
bdf84001
6843b570
8d9a69c5
f002b292
b2890140
4604b08a
f8d3b199
f5b00080
d0074f80
4f00f5b0
f5b0d006
d1055f00
e002211c
e000211d
60a9211e
92016c1a
f402e0e0
b2896180
685bb139
6201210a
f0026e5a
93020301
f402e017
b2895180
685ab141
6201210c
30a8f8d2
0201f003
e00a9203
7100f402
b141b289
2109685b
6e1a6201
0301f002
60a99304
f402e094
b2897180
685ab139
62012108
f0036dd3
92050201
f002e7f1
b2b60604
d0312e00
8beab11d
42828a68
7d68d315
68e3b130
4620b11b
47984629
4618e000
b1126962
46294620
69e14790
2500b111
460d83cd
d1012802
4608e0a5
6f1a6863
d5fc0712
686a6919
b11ab2c9
8a6e8beb
d803429e
4016f240
e08a6220
69e154d1
1c538bca
e08283cb
0110f002
2900b289
b11dd042
8a288ba9
d31f4281
b1587d28
b14268a2
46204629
68634790
f0216b19
631a0210
4610e000
b1136923
46294620
69e14798
2500b111
460d838d
d1062801
8a1a6863
01fff022
e0008219
1e434630
d9542b01
b1196829
8a2b8baa
d8074293
8a036860
01fff023
f2408201
e0444317
5c896863
f0228a1a
430a02ff
69e3821a
1c4a8b99
e03a839a
0f01f012
685bd009
6c5a6201
f00260a9
93060301
bb3b69a3
f002e05f
b2810002
2101b131
6221685a
40086c90
e0169007
0008f002
b139b281
2103685a
6cd06221
0301f000
e00a9308
0220f002
b170b290
2105685a
6d106221
0301f000
60a99309
2b0069a3
4620d039
47984629
f240e035
62234312
2801e031
6861d107
2084f891
0301f042
3084f881
2802e027
7d28d125
6863b180
1088f893
0202f041
2088f883
f8937da8
f000208c
f0220107
43080007
008cf883
b1837d6b
f8906860
f0411088
f8800201
7deb2088
2090f890
0107f003
0307f022
f880430b
b00a3090
b082bd70
1001f04f
4770b002
47702047
d80b2901
f8936843
f0012098
f0220101
43010001
1098f883
47702000
4001f240
68434770
f042881a
80180040
b1a94770
d1162901
2b01b94a
88996843
f441bf0c
f3626180
8099218a
2a01e006
6843d109
f442889a
80985000
47702000
4004f240
f2404770
47704001
47702028
47702028
1181eb00
40106b88
79034770
0101f001
0201f023
71014311
7a034770
0101f001
0201f023
72014311
eb004770
f8911181
f0433028
f8810001
47700028
1181eb00
3028f891
0001f023
0028f881
eb004770
f8911181
f043302c
f8810001
4770002c
1181eb00
302cf891
0001f023
002cf881
eb004770
6bcb1181
0202ea23
477063ca
1181eb00
431a6bcb
477063ca
1282eb00
40086b90
68434770
f0017c18
f0200103
ea400018
741901c1
f0027c18
f0200207
430a0107
4770741a
d80a2903
f001e8df
08060402
47706082
477060c2
47706102
47706142
d80a2903
f001e8df
08060402
47706082
477060c2
47706102
47706142
6984b5f8
f8946842
eb02102f
46051181
07f06b8e
6a2bd54a
428369a0
69e0d202
d3034283
5206f240
e03f84aa
0032f894
28013801
6a08d80d
f8216921
f8940013
eb02002f
6a481180
f8216961
33010013
f894622b
1ec10032
d8182901
302ff894
1083eb02
6a016923
0017f3c1
f8436a29
f8940021
6963002f
1280eb02
6a2a6a51
0017f3c1
0022f843
1c486a29
6a2b6228
429369a2
69e1d202
d307428b
b12b68ab
46214628
f44f4798
84a060a1
d55b06f1
102df894
d1572901
68a069eb
d2024283
429368e2
2300d301
f894e04c
1e481031
d8182801
f894686a
6827102f
1181eb02
7013f837
f3676a08
62080017
702ff894
eb026861
f8311287
6a510013
f3603301
62510117
f89461eb
1ec20031
d8192a01
f894686a
69eb102f
eb026827
f8571181
6a087023
0017f367
f8946208
6861702f
1287eb02
0023f851
33016a51
0117f360
61eb6251
68a269e8
d2024290
428868e1
68ebd30a
4628b133
47984621
5007f240
e00184a0
302df884
d50e07b2
5206f240
f89484aa
6869302f
01821c58
68e9588b
696bb119
46214628
06b34798
f240d50f
84a85005
202ff894
1c536869
1083eb01
684368e9
692ab119
46214628
bdf84790
6984b5f8
f8946843
eb03202f
46051182
07b26b8e
f240d50b
84825206
102ff894
01911c4a
68c3585b
4621b10b
06f14798
f894d55a
2801002d
69ebd156
429368a2
68e1d202
d301428b
e04b2300
0031f894
2a011e42
686ad818
102ff894
eb026827
f8371181
6a087013
0017f367
f8946208
6861702f
1287eb02
0013f831
33016a51
0117f360
61eb6251
0031f894
2a011ec2
686ad819
102ff894
682769eb
1181eb02
7023f857
f3676a08
62080017
702ff894
eb026861
f8511287
6a510023
f3603301
62510117
69e861eb
429068a2
68e1d202
d3094288
b12b68eb
46214628
20004798
e00161e8
302df884
d54907f2
69a16a2b
d202428b
429369e2
f240d303
84ab5306
f894e03e
38010032
d8132801
702ff894
c004f8d5
1087eb0c
69206a07
7013f820
702ff894
1087eb0c
69606a47
7013f820
622b3301
0032f894
2b011ec3
f894d814
f8d5702f
6a2bc004
1087eb0c
69206a07
7013f820
702ff894
1087eb0c
69606a47
7013f820
622b3301
42886a28
4290d201
68aad306
4621b122
47904628
62292100
d50e06b3
5005f240
f89484a8
6869202f
eb011c53
68ea1083
b1126843
46214628
bdf84790
f0437b03
73010101
00004770
6843b538
781a460c
46054949
f042428b
70180001
4a47d103
60106810
4a46e008
d1054293
5080f502
f36f69c1
61c1314d
29017a61
4a3ed13c
d11c4293
28017860
4b3ed10a
68197922
00527960
0101f041
0080ea42
60194301
2b0178a3
4b37d128
681a79a0
0101f042
00527922
0080ea42
60194301
4830e01c
d1194283
2b017863
7961d109
00887922
0342ea40
0101f043
f7fb482b
78a2fb4f
d1092a01
792079a1
ea43008b
f0420240
48250101
fb42f7fb
78e2686b
eb037960
f0001282
f8920007
f0211034
43010107
1034f882
79a078e2
1282eb03
0007f000
1030f892
0107f021
f8824301
79e01030
d9022807
2a077a22
78e1d81a
1281eb03
010ff000
004cf892
000ff020
f8824301
78e2104c
eb037a20
f0001382
f893010f
f0222048
4308000f
0048f883
bd382000
5001f240
bf00bd38
47050000
46008044
24040400
46008034
24041400
6843b538
781a460c
4605494a
f042428b
70180001
4848d105
f4416801
60020200
4a46e008
d1054293
5080f502
f44169c1
61c25200
28017a60
493ed13c
d11c428b
28017860
4b3ed10a
68197922
00527960
0101f041
0080ea42
60194301
2b0178a3
4b37d128
681a79a0
0101f042
00527922
0080ea42
60194301
4a30e01c
d1194293
2b017863
7961d109
008a7920
0340ea42
0101f043
f7fb482b
78a0faab
d1092801
792279a1
008b4827
0242ea43
0101f042
fa9ef7fb
78e2686b
eb037960
f0001282
f8920007
f0211034
43010107
1034f882
79a078e2
1282eb03
0007f000
1030f892
0107f021
f8824301
79e01030
d9022807
2a077a22
78e1d81a
1281eb03
010ff000
004cf892
000ff020
f8824301
78e2104c
eb037a20
f0001382
f893010f
f0222048
4308000f
0048f883
bd382000
5001f240
bf00bd38
47050000
46008044
24040400
46008034
24041400
460db538
0103f010
d10c4604
f0042228
6868f807
6060682b
78026023
0101f022
46207001
2000bd38
b538bd38
f010460d
46040103
2228d10c
fff2f003
682b6868
60236060
f0227802
70010101
bd384620
bd382000
4605b538
2900460c
80aef000
202ff891
f2002a01
698b80a9
69c8b90b
f894b348
b929102c
2b006923
6960d059
d0562800
494f686b
d10e428b
d1062a01
1028f893
0201f021
2028f883
f893e005
f0222068
f8830001
79180068
0101f040
f8947119
eb03202f
f8931382
f0400028
f8830101
6a231028
d50203d9
2a0068aa
041ad02f
68ebd505
d02a2b00
46214628
6a204798
d50403c3
b11268aa
46214628
4a354790
68136a21
bf4c0448
4380f443
4380f423
68a16013
220061ac
5004f240
84a02301
622a84aa
f88461ea
b909302d
b1f868e0
202cf894
6823b93a
6861b10b
f240b919
84a15101
6868e042
42904a21
f894d110
2b01302f
f890d106
f023302c
f8800101
e005102c
106cf890
0201f021
206cf880
302ff894
6aa26868
1183eb00
f89463ca
b98b302c
202ff894
1382eb00
102cf893
0201f041
202cf883
f0437a03
72010101
f0427b02
73030301
07c16a20
8ca0d402
e00bb281
f2408ca1
b20a5304
d1f6429a
f7ff4628
e7f5fc2d
5101f240
bd38b208
47050000
46008068
4605b538
2900460c
809ef000
202ff891
f2002a01
698b8099
69c8b90b
f894b348
b929102c
2b006923
6960d04d
d04a2800
4947686b
d10e428b
d1062a01
1028f893
0201f021
2028f883
f893e005
f0222068
f8830001
79180068
0101f040
f8947119
eb03202f
f8931382
f0400028
f8830101
6a231028
d50103d9
b32268aa
d504041a
b30368eb
46214628
6a204798
d50403c3
b11268aa
46214628
68a24790
230061ac
5104f240
84a12001
622b84ab
f88461eb
b90a002d
b1f968e1
302cf894
6820b93b
6862b108
f240b91a
84a05001
6869e03e
42994b1f
f894d110
2801002f
f891d106
f020002c
f8810201
e005202c
206cf891
0301f022
306cf881
102ff894
6aa0686b
1281eb03
f89463d0
b969102c
002ff894
1280eb03
102cf892
0001f041
002cf882
f0427a1a
72190101
07d86a23
8ca3d402
e00bb298
f2408ca0
b2025104
d1f6428a
f7ff4628
e7f5fc59
5001f240
bd38b200
47050000
4801b082
4770b002
00010201
4770203b
f0437d03
75010101
7e034770
0101f043
47707601
1181eb00
3050f891
0001f043
0050f881
eb004770
f8911181
f0433054
f8810001
47700054
29034770
e8dfd820
0902f001
f8901810
f0433034
f8800102
e00c1034
110cf890
0202f041
210cf880
f890e005
f0422124
f8800302
20003124
f8904770
f043313c
f8800102
e7f6113c
7001f240
29034770
e8dfd820
0902f001
f8901810
f0233034
f8800102
e00c1034
110cf890
0202f021
210cf880
f890e005
f0222124
f8800302
20003124
f8904770
f023313c
f8800102
e7f6113c
7001f240
b5104770
d82f2903
f001e8df
25100702
85838d81
85028d03
f8b0e01b
f8a01104
f8b03104
f8a03100
e0122100
111cf890
0301f003
0401f021
f8804323
f890311c
f0021118
f0210201
ea440401
f8800302
20003118
f8b0bd10
f8a01134
f8b03134
f8a03130
e7f42130
7001f240
2903bd10
e8dfd80e
0402f001
6bc00a07
f8d04770
47700114
012cf8d0
f8d04770
47700144
7001f240
29034770
e8dfd80e
0402f001
6b800a07
f8d04770
47700110
0128f8d0
f8d04770
47700140
7001f240
29014770
0049d802
10f0f8c0
f0037913
f8900103
f0233148
ea430306
f8800141
78131148
010ff003
30f8f890
030ff023
f880430b
885230f8
20fcf8c0
b5304770
2b01780b
f240d902
bd307004
d8692a03
f002e8df
35351802
784cb95b
d8f22c03
030ff004
4080f890
040ff024
f8804323
780b3080
d1382b01
2b03788b
f003d8e3
e016030f
784cb963
d8dc2c03
f89000a3
f0034080
f024030c
4323040f
3080f880
2b01780b
788bd121
d8cc2b03
f004009c
f890030c
f0244084
4323040f
b943e013
2c03784c
f890d8bf
f0233080
f880040f
780b4080
d1082b01
2c03788c
f890d8b3
f0233084
f880030f
780b3084
f102b95b
78cd0311
4033f810
053ff005
043ff024
f800432c
780b4033
d10e2b01
eb003211
790900c2
f0017903
f023023f
4311013f
e0027101
7001f240
2000bd30
2903bd30
e8dfd820
0902f001
f8901810
f0433034
f8800104
e00c1034
110cf890
0204f041
210cf880
f890e005
f0422124
f8800304
20003124
f8904770
f043313c
f8800104
e7f6113c
7001f240
29034770
e8dfd820
0902f001
f8901810
f0433034
f8800101
e00c1034
110cf890
0201f041
210cf880
f890e005
f0422124
f8800301
20003124
f8904770
f043313c
f8800101
e7f6113c
7001f240
67c14770
67814770
60c14770
68434770
60414319
68834770
60814319
68004770
47704008
d81a2a03
f002e8df
130c0602
43116b02
e00a6301
3108f8d0
f8c04319
e0041108
2120f8d0
f8c04311
20001120
f8d04770
43193138
1138f8c0
f240e7f7
47707001
d8022a03
20006501
f2404770
47707001
d8022a03
20006541
f2404770
47707001
d8062907
fa032301
f8c0f101
200010d0
f2404770
47707004
d8062907
fa032301
f8c0f101
200010d4
f2404770
47707004
10c8f8c0
f8c04770
477010cc
d8052907
f101fa02
10d8f8c0
47702000
7004f240
29074770
fa02d805
f8c0f101
200010dc
f2404770
47707004
10e0f8c0
f8c04770
477010e4
d8082907
30e8f8d0
f101fa02
f8c04319
200010e8
f2404770
47707004
d8082907
30ecf8d0
f101fa02
f8c04319
200010ec
f2404770
47707004
f8c02301
477030f0
f8c02301
477030f4
47706781
477067c1
d8062a03
f8303216
f8203022
20001022
f2404770
47707004
3148f890
0101f001
0208f023
01c1ea42
1148f880
f8904770
f0013148
f0230101
43110201
1148f880
2a034770
e8dfd82a
0a02f002
8e031f14
0207f001
0107f023
8602430a
f8b0e012
f0013108
f0230107
43110207
1108f8a0
f8b0e008
f0013120
f0230207
430a0107
2120f8a0
47702000
3138f8b0
0107f001
0207f023
f8a04311
e7f31138
7001f240
2a034770
e8dfd80e
0402f002
03090b06
0349e002
0389e000
10e0f8c0
47702000
e7f903c9
7001f240
f8c04770
f8c020e0
477010e0
680bb538
460d6804
d0332b00
d50107e2
47982000
d50207a0
20016829
07614788
682ad502
47902002
d5020722
2003682b
06e34798
6829d502
47882004
d50206a0
2005682a
06614790
682bd502
47982006
d5020622
20076829
05e34788
682ad502
47902008
7000f414
2009d006
4798682b
bd382000
7004f240
b082bd38
2002f04f
4770b002
23082000
0003f363
f3612102
47701005
d8092901
b9117803
0101f043
f043e001
70010102
47702000
4001f241
23004770
47706003
2300b510
d2044293
f8416844
33044023
bd10e7f8
47706001
47706041
43196d03
47706501
43196d43
6d816541
6582430a
6ec34770
66c14319
430a6f01
47706702
43196e03
6e416601
6642430a
6f834770
67814319
430a6fc1
477067c2
3084f8d0
f8c04319
f8d01084
430a1088
2088f8c0
f8d04770
43193090
1090f8c0
1094f8d0
f8c0430a
47702094
30a8f8d0
f8c04319
f8d010a8
430a10ac
20acf8c0
f8d04770
4319309c
109cf8c0
10a0f8d0
f8c0430a
477020a0
43196e83
47706681
43196dc3
477065c1
43196f43
47706741
3080f8d0
f8c04319
47701080
308cf8d0
f8c04319
4770108c
3098f8d0
f8c04319
47701098
30a4f8d0
f8c04319
477010a4
d9012903
d80f2a03
f0017e03
f023010f
4319030f
7f037601
020ff002
010ff023
7702430a
47702000
1002f640
6a434770
62414319
68034770
d402061a
02136802
69c2d503
61c14011
69834770
61814019
6a834770
62814319
00004770
f04f4b03
601a32ff
43116902
47706101
46110010
431968c3
477060c1
43196943
47706141
40086880
b9114770
b2886a01
29014770
6a00d102
47700c00
1001f640
b9114770
b2886a41
29014770
6a40d102
47700c00
1001f640
b91a4770
f3616a83
e0040343
d1032a01
f3616a83
62834353
f8d04770
401930b0
10b0f8c0
b1094770
d1002901
47706001
6f42b919
0140f042
2901e004
6f43d103
0100f443
47706741
d8042901
0300f04f
6001d105
f640e004
b2001002
60034770
e7fa4618
d8032901
2202b931
e0016002
1101f640
4770b208
3300f44f
21006003
2901e7f8
b931d803
60022208
f640e001
b2081101
f44f4770
60032300
e7f82100
d8052901
b9396a83
0201f043
e0016282
1101f640
4770b208
3180f443
21006281
2a01e7f8
6bc3d805
f361b93a
63c3230f
f640e001
b2101201
f3614770
63c3631f
e7f82200
d80c2a01
b919b98a
f3636a82
e004224b
d1072901
f3636a82
62821288
f640e002
e0001101
b2082100
b9214770
f3636a82
6282625b
2901e7f7
6a82d1f4
5298f363
2a01e7eb
b98ad80c
6bc2b919
0202f363
2901e004
6bc2d107
02c5f363
e00263c2
1101f640
2100e000
4770b208
6bc2b921
4212f363
e7f763c2
d1f42901
f3636bc2
e7eb42d5
b5702901
460e4604
d83b461d
d13d2900
6ae38898
030ff360
88e962e3
f3616ae0
62e0401f
f0136aa3
d1030f0e
f4116aa1
d0012f60
63606968
d1172a01
06c16aa0
682bd508
f640b913
e01d1602
46292009
47984632
f4126aa2
d02c1380
2b00682b
200ad0f1
46324629
e0244798
6ba2b9ce
f36089a8
63a2421f
6c2389e9
030ff361
e0016423
1601f640
bd70b230
6b038919
030ff361
89686303
f3606b21
6321411f
6ba6e7c0
f3628a2a
63a6060f
6c238a69
431ff361
26006423
b510e7e6
8894b951
f3646ac3
62c3030f
6ac188d2
411ff362
e00b62c1
d10b2901
6b038911
030ff361
89526303
f3626b01
6301411f
e0012000
1001f640
bd10b200
4613b570
b981460c
f0116881
d0020508
20046815
6880e01c
0004f010
6814d02a
20034611
47a0462a
2901e015
6885d108
2500f415
6882d10a
2280f412
e010d00b
d1142902
f4126882
d0062500
2008681d
46224619
230047a8
6881e00d
2080f411
681ed008
46192007
47b04622
f640e7f3
e0001301
b2184603
b082bd70
3081f44f
4770b002
20002304
0002f363
f3612108
220200c6
10caf362
f3632326
f44020d0
47703000
4770203c
60832301
23004770
47706083
d8052901
f3616803
60031386
47702000
2001f241
29014770
6803d805
13c7f361
20006003
f2414770
47702001
f3616803
60035356
47702000
f3616803
60031305
47702000
f3616803
60032309
47702000
47706101
61032300
6a804770
62c14770
6b004770
6b404770
b0824770
93016c83
b0029801
b5704770
0383eb01
42942400
b2a0d101
6805bd70
2e006a2e
f833d0f9
f8b51024
f8a56060
34011060
b570e7ef
0383eb01
42942400
b2a0d101
6805bd70
2e016a6e
6e29d0f9
f843b289
34011024
b5f0e7f1
0343eb01
42942400
d00ab2a6
6a2f6805
f833b93f
f8b51014
f8a56060
34011060
4630e7f1
b530bdf0
0343eb01
42942400
6805d008
29006a69
6e29d0fc
1014f823
e7f43401
bd30b2a0
2400b5f0
b2e64294
4630d101
6805bdf0
2f006a2f
18ced1f9
7060f8b5
34015d36
6060f8a5
b570e7ee
42942400
6805d008
2e006a6e
6e2ed0fc
552e18cd
e7f43401
bd70b2e0
f8802300
f8803035
47703036
6a826a43
b5106859
fbb16854
f013f3f4
d1010f01
e0046094
fbb14c04
4361f1f3
68006091
8a81b29a
bd108282
000f4240
f010b510
d16d0403
2b00684b
680ad06c
e8806241
6094000c
68036a42
29017ad1
681ad803
1286f361
6a41601a
7a896803
d8032901
f361681a
601a12c7
6a416803
7a09681a
5256f361
6803601a
681a6a41
f3617b09
601a1205
68036a41
f0027b8a
7e1a010f
020ff022
761a430a
68036a41
f0027c0a
7f1a010f
020ff022
771a430a
68036a41
f0027c8a
f8930101
f022204c
ea420202
f8830141
6803104c
7d116a42
204cf893
0101f001
0201f022
f883430a
6a41204c
7d8a6803
010ff002
2050f893
020ff022
f883430a
6a412050
7e0a6803
010ff002
2054f893
020ff022
f883430a
bd102054
bd102000
bd104618
d80a2903
f001e8df
08060402
47706082
477060c2
47706102
47706142
b1104b05
7080f44f
681ae002
7080f422
20006018
bf004770
46008014
6ac6b5f8
429e684b
460d4604
6987d206
22016809
47b84633
62e01980
68696ae2
d30c428a
b15368e3
26004805
68e262c6
46294620
f8844790
f8846035
bdf86036
44020000
68cab570
42956b05
d3064604
b15b6903
4a064798
62d12100
69c6bd70
22016889
47b0462b
63201940
bf00bd70
44020000
6803b538
6b196a05
460407cb
f890d508
2a012035
682bd104
4629b113
ffb6f7ff
7a416a60
d1032902
f2416823
661a2234
6b216a20
429968c3
6882d205
4620b11a
f7ff4629
6a20ffc5
68436ae1
d30e4299
49076822
f8842000
61100035
68a362c8
46294620
6a204798
2204f241
bd386142
44020000
460db538
b9104604
2001f241
2900bd38
62a1d0fa
1e59784b
d8f5291f
2a00686a
f7ffd0f2
6820fecf
68026a63
f3617a59
60022209
68236aa0
29107841
1e48d901
681ae007
4214f36f
6aa0601a
78416823
681a1e48
4214f360
78a9601a
1e486823
8899b282
6aa1809a
780a6823
4b0b611a
62d82000
22016821
786b608a
d9032b10
4a084907
e00761a1
4b07d003
61a34a07
4907e002
61a14a07
bd3861e2
44020000
0030cd37
0030cd5f
0030cdcd
0030cdf3
0030cd83
0030cdab
460cb538
28004605
2900d033
7e0bd031
d9032b0f
2001f241
bd386148
2202f241
62292300
2201614a
3034f880
2035f880
3036f880
62c36303
009b690b
68c2d501
69204790
d50300c2
4628692b
47984621
21054a09
692062d1
db012800
bd382000
f7ff4628
6963ff37
2102f241
d0f7428b
f241e7f4
bd382001
44020000
4770203c
60832301
23004770
47706083
d8052901
f3616803
60031386
47702000
2001f241
29014770
6803d805
13c7f361
20006003
f2414770
47702001
d8052902
f3616803
60035356
47702000
2001f241
29024770
6803d805
1305f361
20006003
f2414770
47702001
d8052904
f3616803
60032309
47702000
2001f241
6a804770
62c14770
6b004770
6b404770
6c804770
23004770
3038f880
3039f880
b5704770
0383eb01
20004605
d00a4290
6a26682c
f833b13e
f8b41020
f8a46060
30011060
bd70e7f2
eb01b570
46050383
42902000
682cd009
2e016a66
6e21d005
f843b289
30011020
bd70e7f3
eb01b5f0
24000343
b2a64294
6805d00a
b93f6a2f
1014f833
6060f8b5
1060f8a5
e7f13401
bdf04630
eb01b530
24000343
d0054294
6e296805
1014f823
e7f73401
bd30b2a0
2400b5f0
b2e64294
4630d101
6805bdf0
2f006a2f
18ced1f9
7060f8b5
34015d36
6060f8a5
b5f0e7ee
42942400
d101b2e6
bdf04630
6a6f6805
d0f92f01
18cd6e2e
3401552e
f010e7f1
d1780203
6241680b
609a6003
68036a41
290179c9
681ad803
1286f361
6a41601a
79896803
d8032901
f361681a
601a12c7
68036a41
29027909
681ad803
5256f361
6a41601a
7a096803
d8032902
f361681a
601a1205
7a596a43
681a6803
f442b111
e0016280
228af361
6a41601a
7a8a6803
010ff002
f0227e1a
430a020f
6a41761a
7b0a6803
010ff002
f0227f1a
430a020f
6a41771a
7c8a6803
010ff002
2050f893
020ff022
f883430a
6a412050
7d0a6803
010ff002
2054f893
020ff022
f883430a
6a412054
7c0a6803
0101f002
204cf893
0201f022
f883430a
6a41204c
7b8a6803
0101f002
204cf893
0202f022
0141ea42
104cf883
20004770
29034770
e8dfd80a
0402f001
60820806
60c24770
61024770
61424770
00004770
41f0e92d
f015690d
46045300
d0084688
22026803
68c364da
d0312b00
e8bd4798
f01581f0
6ac66580
d00f684a
d3054296
3038f880
3039f880
81f0e8bd
69854911
47a82201
62e11981
81f0e8bd
d3024296
62dd4b0d
2201e010
68094633
47b86987
3004f8d8
42981980
d30962e0
62cd4906
f2416a20
82822204
5038f884
5039f884
81f0e8bd
00300ba0
45010000
690bb5f8
5380f013
460d4604
6803d005
64da2201
b9cb6903
6b06e019
429668ca
f241d306
63422204
48096c82
bdf862c3
69c76889
46332201
68e947b8
42881980
d3046320
b1136923
46294620
bdf84798
45010000
6803b538
6b196a05
460407cb
f890d508
2a012038
682bd104
4629b113
ff80f7ff
6b216a20
429168c2
6883d205
4620b11b
f7ff4629
6a20ffbb
68426ae1
d3084291
23004808
3038f884
6a2162c3
2204f241
6a23828a
68d96b20
bf244288
2105f241
bd388299
45010000
2800b510
2900d02f
6a42d02d
79546281
2c046803
681ad803
2209f364
6a83601a
6803785c
2c10681a
34fff104
f364bf8c
f3644214
601a0203
23006802
62c32401
78496094
d9032910
61814908
e0074908
4a08d003
61824908
4a08e002
61824908
461861c1
f241bd10
bd102001
0030d22b
0030d251
0030d2b9
0030d2df
0030d275
0030d29d
460db538
28004604
2900d02f
7d8bd02d
d82a2b0f
2202f241
62212300
2201828a
2038f880
3039f880
63036343
690b62c3
d501009b
479068c2
00c26928
6923d503
46294620
4a0a4798
62d12105
28006928
2000db01
4620bd38
ff5cf7ff
1014f9b5
2302f241
d0f64299
f241e7f3
bd382001
45010000
47706001
b2c06800
68034770
611a2220
68034770
611a2200
68034770
4311685a
47706059
685a6803
60594011
68034770
47706998
61196803
68034770
47706958
10fff240
b5384770
68ac6805
0307f004
d1052b07
69c36feb
d0422b00
e02c210c
0206f004
d1222a06
f013696b
d0030402
b3b369c3
e0202107
0204f013
69c3d003
2108b37b
f013e02b
d0030408
b34369c3
e0252109
0210f013
69c3d003
210ab30b
061be01d
69c3d51d
210bb1db
f014e018
69c30202
b1a3d003
22002101
f004e010
290c010c
b163d102
e0092106
0404f014
b133d002
e0032102
b113692a
46222103
bd384798
477068c0
47706980
61c1b111
47702000
6001f240
68034770
2040f893
0002f042
0040f883
47702000
f8936803
f0222040
f8830002
20000040
b5084770
22042100
fba4f002
bd082000
460fb5f8
28004606
4b22d040
5196f5a1
d83b4299
f0014610
4604fd31
460d4638
fd2cf001
4b1c2200
fd9ef001
460b4602
46294620
fec2f001
4604460d
ffa6f001
60f12180
20c0f896
073ff022
70c0f886
2700b280
b2c36037
60f76077
0a0160f1
60716033
fd1af001
460b4602
46294620
fbc6f001
4b092200
fd76f001
ff86f001
f8c6b280
60f700c0
bdf84638
6001f240
bf00bdf8
008c8d40
40300000
40500000
41f0e92d
4605780a
b2c41f50
460b2c04
492cd805
5d0e190f
8005f897
f04fe002
26030800
7c5c795a
28011e50
f046bf98
2c000604
240fbf14
60ac2407
29027999
2903d006
2901d007
f044d107
e0040410
0420f044
f044e001
79df0430
d0062f02
d0072f03
d1072f01
0440f044
f044e004
e0010480
04c0f044
7b187b5a
bf142a00
27002720
2f00b118
2730bf14
7b992710
7bdab131
f046b912
e0010608
0618f046
46286899
f44fb909
695a31e1
ff58f7ff
431f692b
60ac612f
f8c560ee
e8bd80cc
bf0081f0
00300bf8
41f0e92d
2058f890
f0424604
f8840001
460b0058
b1297909
5058f894
0602f045
6058f884
1f7a781f
2804b2d0
493cd805
7aae180d
800ff895
f04fe002
26030800
b98778df
2040f894
0001f042
0040f884
f8947919
29015040
f025bf0c
f0450502
f8840502
789f5040
f894b12f
f0422058
f8840010
f8940058
f0411058
f8840520
795f5058
79997c58
2a011e7a
f046bf98
28010604
2509bf0c
29022501
2903d006
2901d007
f045d107
e0040510
0520f045
f045e001
79df0530
d0062f02
d0072f03
d1072f01
0540f045
f045e004
e0010580
05c0f045
7b187b5a
bf142a00
27002720
2f00b118
2730bf14
7b992710
7bdab131
f046b912
e0010608
0618f046
46206899
f44fb909
695a31e1
fec6f7ff
431f6923
60a56127
f8c460e6
e8bd80cc
bf0081f0
00300bf8
460db570
46064614
2100b168
f0022220
6035fa53
46287863
b1134621
ff5ef7ff
f7ffe001
4630fef7
b530bd70
b1aab1b1
68042300
07ed68a5
6fe5d40b
d5f907ad
602556cd
330168c4
42933401
d1f060c4
6fe5e006
0f02f015
e001d1ef
6301f240
bd304618
4607b5f8
460e4615
b152b159
46312400
4638462a
ffd7f7ff
44041a2d
d1f64406
f240e001
46206401
b530bdf8
b172b179
68042300
f0156965
d00a0f01
54cc6824
33016984
42933401
d1f26184
f240e001
46186301
b5f8bd30
46154607
b159460e
2400b152
462a4631
f7ff4638
1a2dffde
44064404
e001d1f6
6401f240
bdf84620
f8d36803
07d220cc
f893d50b
f04000cc
f8830202
f89320cc
f88320c4
200010c4
f44f4770
47707081
47f0e92d
46062902
46984691
a020f8dd
68446807
69f8d002
e0052161
33fff102
d9052b01
215b69f8
f04f6041
e05035ff
69f86882
30086851
7b304788
25004623
da384285
f203461c
78616314
f240bb89
46206214
f9aaf002
0920f049
70622201
9002f884
0f00f1ba
f8c4d002
e003a60c
f0617ee1
76e0007f
0f01f018
7ee3d003
0201f043
f01876e2
d00d0f04
f3c87ee1
f04103c3
76e00004
2204b90b
b2dae000
2609f884
2608f884
18c3f3c8
860af884
3501e001
7b31e7c4
69f868b3
428d689a
0008f100
4790db04
21176835
e7ab69e8
46284790
87f0e8bd
2400b513
f7ff9400
bd1cff8f
4ff0e92d
1e0eb093
92044604
e8904699
db1a0120
429e7b03
f240dc17
fb076714
eb08fb06
f89a0a0b
f0011002
2a01020f
69ebd005
605a225b
30fff04f
f89ae0b8
93023001
2b013b03
69ebd902
e7f22209
2018f89a
d0022a01
221669eb
f89ae7eb
f89ac019
459c301a
69ebd102
e7e22269
2b049b02
f89ad118
f8da301b
0909660c
f0039600
f7ff0301
b2c6ff49
2800b270
7b21dbd2
dccf4288
8700fb07
3004f8ba
763a2202
e00080bb
68a1b2f6
684f69e8
47b83008
462069e9
f0003150
4607fd80
68a3b948
689969e8
47883008
f06f6820
69c30203
f818e7af
7538000b
0115f107
f8ba4620
f0012004
69eaf90e
6058f882
206c68a3
46396a1a
46834790
d1472800
29009904
f8d9d038
28000000
b273d034
6214f240
8103fb02
091a788b
d10e2a02
88c9688b
201cf8ad
93082810
101ef8ad
2210d902
2000f8c9
a9079804
2a03e018
88cbd11a
202cf8ad
0208f101
302ef8ad
f101920d
f101030c
31140210
930e281c
9110920f
201cd902
0000f8c9
a90b9804
2000f8d9
f806f002
f240b270
fb036314
f89a8100
2204001a
704a1c43
301af88a
463a69e9
46203150
fd2af000
69e868a1
3008688a
f1bb4790
f47f0f00
b270af45
e8bdb013
e92d8ff0
46984ff0
f240b08f
f8d06314
9201b004
fa01fb03
46042900
68054689
070aeb0b
7b02db05
dc024291
28047878
69ebd002
e0222109
69e868a1
3008684e
7ba347b0
d0042b01
f8c79a01
f8c78604
f8d72600
b11005fc
29017ba1
69e9d043
31504620
fcd1f000
b9504606
69e868a1
3008688a
68204790
f06f69c3
60590103
2100e02e
f1002207
f0020014
f81bf843
f240300a
459052b4
4690bfa8
46207533
0115f106
f0014642
4620f85d
0119f106
2610f8b7
f84df001
f88069e8
68a19058
6a0b206b
47984631
69e9b170
46204632
f0003150
68a2fcb3
689369e8
47983008
38fff04f
2600e068
2a017ba2
f8d7d121
f8d705fc
454015f8
4680bf38
311c1879
98014642
ff64f001
05fcf8d7
35f8f8d7
bf2c4540
0000ebc8
f8c72000
f8d705fc
eb0315fc
f8c70208
b92125f8
15f8f8c7
f8d7e001
9b198604
d0322b00
68129a1a
d02e2a00
88f978b8
2b020903
68b8d10d
300cf8ad
90042a10
100ef8ad
991ad902
600b2310
a9039819
2003e017
0308f107
001cf8ad
101ef8ad
f1079309
f107010c
f1070010
2a1c0314
900b910a
d902930c
211c9a1a
98196011
9a1aa907
f0016812
69e9ff17
31504620
f0004632
68a3fc47
689969e8
47883008
b00f4640
8ff0e8bd
b086b570
2500ac06
5d04f844
95019e0a
94029600
ff15f7ff
bd70b006
4ff8e92d
0800f1b1
46934604
0420e890
7b03db02
dd024598
220969eb
f240e028
fb036314
eb0af908
787a0709
d00a2a04
28017e38
4638d007
461a2100
ff7cf001
e8bd2000
68a18ff8
684e69e8
47b03008
462069e9
f0003150
4606fbea
68a2b968
689169e8
47883008
69c36820
0203f06f
f04f605a
e8bd30ff
f1bb8ff8
46200f01
0114f106
2200d107
ff75f000
f1064620
88ba0116
f81ae007
f0002009
4620ff6c
0116f106
f0002200
69efff66
8058f887
463168a3
20436a1a
69e94790
31504607
46204632
fbccf000
69e868a1
3008688b
2f004798
f04fbf14
200030ff
8ff8e8bd
4ff8e92d
68466807
69f94689
46053150
469b4692
fb9bf000
28004604
8085f000
0814f100
22892100
f0014640
f240ff15
fb036314
46416609
090278b0
46282a02
2204d105
ff27f000
61e368b3
2206e00e
ff21f000
0308f106
021cf104
0118f106
0b04f853
f842428b
d1f90b04
f1044628
88b20118
ff0ff000
f1044628
88f2011a
ff09f000
f1044628
fa1f0116
f000f28a
f1baff02
46280f02
012cf104
fa1fd10a
f000f28b
f894fef8
f042209b
f8840102
e002109b
f0002200
7ef0feee
d50507c3
3032f894
0201f043
2032f884
101bf996
da052900
009bf894
0301f040
309bf884
f0027ef2
b2c80104
f894b128
f043309b
f8840204
f894209b
f041109b
f8840010
f896009b
f884660a
69fb609c
9058f883
462168aa
20426a16
69f947b0
31504606
46224628
fb2cf000
f04fe001
463036ff
8ff8e8bd
47f0e92d
46041e0f
68436805
7b01db19
dc16428f
6614f240
3607fb06
9002f896
090ff009
0f01f1b9
69ebd006
6058205b
30fff04f
87f0e8bd
a001f896
0f02f1ba
69ebd002
e7f22009
800ff890
bfa84542
68824690
685369e8
47983008
46204639
46434652
ff32f7ff
b9284607
70702003
9018f886
8019f886
69e868a1
3008688a
2f004790
f04fbf14
200030ff
87f0e8bd
41f0e92d
0800f1b1
46074615
68426806
7b01db08
dc054588
6414f240
2408fb04
b9107860
230969f0
b915e012
230e69f0
882ae00e
d1012a02
e0022b10
d1012a03
d1032b1c
ebb278a3
d0061f13
236169f0
f04f6043
e8bd30ff
68b981f0
684a69f0
47903008
28028828
686bd102
e00b60a3
0308f105
0208f104
0118f105
0b04f853
f842428b
d1f90b04
886d78a2
010ff002
80e52901
2200d104
46414638
e0084613
d10a2902
28017860
4638d107
22044641
f7ff2300
4605fec3
2304b910
25007063
69f068ba
30086891
2d004788
f04fbf14
200030ff
81f0e8bd
43f8e92d
0800f1b1
46174604
0220e890
7b02db09
dc064590
6614f240
9608fb06
28017870
69e9d002
e0312209
b913b107
220e69e9
8839e02c
d1012902
e0022b10
d1012903
d1032b1c
ebb178b3
d0021f13
226169e9
68a2e01c
685169e8
47883008
88792300
461a7b20
3201e001
4282b2d2
eb09d013
f2030703
88bf6314
d1f4428f
69e868a1
3008688b
68204798
226269c1
f04f604a
e8bd30ff
78b783f8
f00780b1
2802000f
2204d109
46414620
f7ff2300
2204fe59
70724607
2302e002
27007073
69e868a1
3008688b
2f004798
f04fbf14
200030ff
83f8e8bd
2300b530
7b026844
42904618
5ce5da06
f203428d
d0036314
e7f63001
30fff04f
b510bd30
7b026843
42902000
889cda09
d102428c
2c017e1c
3001d005
6314f203
f04fe7f3
bd1030ff
e92d29ef
460741f0
0048e890
2500d10f
429d7b3b
4630da09
f2402100
f0016214
3501fd3d
6614f206
e8bde7f2
29ee81f0
6514f240
69dcd11f
2058f894
6502fb05
f8b54634
25008004
429d7b3b
88a0da11
d10a4540
f00178a1
2a01020f
4620d105
f2402100
f0016214
3501fd19
6414f204
e8bde7ea
fb0581f0
7e236401
d1072b01
b1bb7ea3
1e592003
76a17060
81f0e8bd
d1082b02
f7ff88a1
b2c0ffa0
6600fb05
1e4a7eb1
462076b2
462a2100
41f0e8bd
bcf4f001
81f0e8bd
030ff001
2b010909
202cbf14
29032038
3014bf08
7382f5c0
4282b298
1a12d90b
2001b292
f5b21c41
b2c87f00
f5a2d904
b29a7300
2001e7f6
f0014770
0909000f
bf142801
2338232c
bf082903
f5c33314
2a017082
d003b280
eb003a01
b2982342
e92d4770
469b4ff8
68066843
6414f240
46052900
4692460f
3401fb04
7b00db02
dd024281
210969f0
78a3e008
020ff003
d1072a02
b9507860
215b69f0
f04f6041
e09539ff
d1022a01
29047861
9a0bd1f4
ebb18811
d0021f13
210e69f0
6a33e7ee
68aa980d
69f06198
30086851
78a34788
000ff003
d1122802
2a047862
4628d00f
22044639
f7ff2300
4681fd51
68aab128
689369f0
47983008
2104e06a
f8947061
f0088002
2b02030f
2b01d010
7ee0d111
d41107c1
0202f000
f240b2d3
f24051aa
2b0050b4
4602bf0c
e007460a
62b8f44f
f240e004
e00152b4
526ef240
f0037ee3
b2c80104
bfb8455a
b3604693
9609f894
0f00f1b9
6829d109
69c868ab
22696899
69f06042
47883008
4628e799
fa1f4641
f7fff28b
4548ff45
4628d906
464a4641
ff5bf7ff
e0064683
d9044581
0c09ebc0
c609f884
2200e002
2609f884
69f49b0d
21abb913
69f4e001
68a821ff
465a7321
9b0b6a44
46384651
68aa47a0
69f04604
30086893
2c004798
46d9bf0c
39fff04f
e8bd4648
e92d8ff8
684447f0
6514f240
4401fb05
78a6b090
8060f8dd
c064f8dd
093688e5
46862e02
4692460f
d10e4699
f8ad68a4
94066014
9401ac05
f8ad2410
f8cd5016
94028000
c00cf8cd
2303e01c
5026f8ad
3024f8ad
0508f104
3418a80b
68694606
c6036828
42a53508
d1f74630
221ca909
92029101
8000f8cd
c00cf8cd
46394670
464b4652
ff03f7ff
e8bdb010
b51387f0
94009c04
94012400
ffb3f7ff
b51fbd1c
94009c06
94019c07
94029c08
94032400
feedf7ff
bd10b004
9d06b5f8
4608461f
4616460c
22082100
fba2f001
f2f5fbb7
00811c50
42ab1a7b
1872d312
21006066
42ab3104
6860d90a
88605042
80603001
30018820
19528020
e7f11b5b
bdf82000
30fff04f
b5f8bdf8
460f6883
69984605
887c4780
68aeb924
479069f2
e0094626
68ab6879
6024f851
3c0169d9
807c2200
47886032
bdf84630
b5706883
4605460c
46166998
88614780
428a8822
68aad105
479869d3
30fff04f
1c4bbd70
6862b299
f8428061
68ab6021
478869d9
bd702000
6883b538
460d4604
47806998
886d68a1
479069ca
bd384628
22044b01
4770601a
4600816c
22044b02
2000601a
bf004770
4600816c
f0002101
0000b954
b5106983
b934681c
20016881
49046aca
46204790
f5a4bd10
38041000
bf00bd10
00300d2c
4e17b5f8
68336801
f0136985
46040702
6880d007
6ac34913
47982002
0001f06f
f7ffbdf8
4601ff88
68a3b940
6ada490e
21014790
f04f7721
bdf830ff
f5021d02
31141000
23106028
f5012002
f44f1100
80ab62c8
81aa60a9
46386030
bf00bdf8
4600816c
00300d5e
00300d8e
4604b538
f7ff6805
4602ffb3
4620b128
0158f105
f93ef000
68a3e004
6ada4906
47902004
f7ff4620
4620ffb5
e8bd2100
f0004038
bf00b8b3
00300dbe
4c0cb510
07516822
f7ffd503
2104ff8f
6821e005
d506078a
ffd4f7ff
4a062102
60116021
6880bd10
6ac34904
47982005
bf00bd10
46008180
41050090
00300df1
31586801
b924f000
784db538
092d6944
6882d107
6ad3490a
47982006
70fff64f
f501e00c
81a31100
60214b06
f5022010
21041200
60a280a0
60192000
bd38b200
00300e13
4600816c
60184b01
bf004770
4600816c
60184b01
bf004770
46008170
f04f4b02
601a32ff
bf004770
4600817c
f04f4b02
601a32ff
bf004770
46008178
60184b01
bf004770
46008178
60184b01
bf004770
4600817c
49034b02
60086018
bf004770
46008180
41050090
460bb508
32fff04f
60192100
7c02605a
d1042a01
68c26880
0008f103
bd084790
6883b538
460d4604
47806998
68a26829
69d3686d
4798400d
bd384628
4604b570
6806460d
ffecf7ff
6829b150
f0004620
3010f867
3020f856
4798b10b
e7fee000
28017c20
68a1d105
0008f105
2100690a
bd704790
b5706883
46046805
460e6998
6b694780
220168a3
f606fa02
636e430e
478869d9
28017c20
68a2d104
003cf105
47986953
b538bd70
46046883
460d6998
68234780
6b5a2101
f505fa01
0505ea22
68a3635d
479069da
b538bd38
46046883
460d6998
68234780
6b9a2101
f505fa01
0505ea22
68a3639d
479069da
b538bd38
46046883
460d6998
68234780
6b9a2101
f505fa01
639d4315
69da68a3
7c204790
d1042801
682068a1
303c694b
bd384798
7c42b510
b2d82300
d2054290
fa042401
3301f403
d0f6420c
7c43bd10
d8074299
31106803
0021f853
f843b910
47702021
47702001
b5086880
68022300
604b600b
814b810b
000cf101
bd084790
6883b5f8
f101460c
4606070c
46386859
47884615
b2828920
6065b912
e0026025
601d6863
89216065
1c4868b3
8122b282
46386899
bdf84788
6883b5f8
f101460c
4605070c
46386859
89264788
b15eb2b6
68268922
68301e53
8121b299
89206020
b90ab282
60626022
463868ab
47886899
bdf84630
b5706883
f101460d
4606040c
46206859
896a4788
b12268b0
46206881
25004788
892de004
46206883
4798b2ad
bd704628
b5706883
050cf101
460e4604
68594628
68a24788
81702001
46286893
bd704798
b5706883
050cf101
460e4604
68594628
68a24788
81702000
46286893
bd704798
4ff7e92d
92016806
69f14689
6843461f
46053150
f7ff9300
4604fd9c
f0002800
f1008098
21000804
f1042210
46400b14
f914f001
221c2100
f0014658
9800f90f
6214f240
f909fb02
0a09eb00
f89a4628
090b1002
46592b02
2204d116
f91df000
68539a0c
46286223
011ef104
f0008852
f89af914
f0000002
2901010f
f04fbf14
f04f0b2c
e0130b38
f0002206
9a0cf906
f1044628
8852011e
f8fff000
0002f89a
010ff000
bf142901
0b40f04f
0b4cf04f
301bf89a
0202f003
b138b2d0
bf8c2f7d
21062108
030beb01
fb83fa1f
f8129a00
75a00009
1003f89a
75e14628
f104b2ba
f0000118
4628f8da
011cf104
f000465a
f104f8d4
f1ab0914
fa19031c
9901f083
301c463a
f001445f
053af807
46414628
f0000d12
7960f8c2
0150f040
71614622
f1064628
f7ff0124
4628fef9
f7ff2101
68abfe79
691a69f0
30102100
69f14790
730e2600
684e4628
31504622
fd1af7ff
f04fe001
463036ff
8ffee8bd
4ff8e92d
f8d0798f
68459000
f101460c
31040a14
f0004606
2f01f8ac
f8d9d10a
0502301c
20006c9b
0d124651
20004798
8ff8e8bd
7da14630
faf0f7ff
f880fa4f
0f00f1b8
b017f894
f04fda03
e8bd30ff
f2408ff8
f1046314
46300118
5508fb03
f887f000
011cf104
46304607
f881f000
7ee84603
d41b0602
c60cf8d5
0f00f1bc
f000d0d5
b2f60602
211cb166
43481e58
f80a18e1
3113b000
560cf8d5
1c7a4640
e7c447a8
464018e1
463a3114
e7be47e0
2a017bb2
f8d5d10d
290015fc
18e1d1c5
001cf105
463a3114
ff78f000
75fcf8c5
f8d5e00c
b1380600
311418e1
f000463a
f8c5ff6d
e0017604
0604f8c5
f00378ab
2802000f
f104d116
4630011e
f839f000
80e878aa
29020911
0320f104
681ad102
e00760aa
34303508
0b04f853
f84542a3
d1f90b04
001cf8d9
296b7b01
af7ff47f
240068b3
695a7304
47903010
7b40e777
b9100a13
704b700a
704a4770
4770700b
7b44b510
0a100c13
7048b92c
700a0e10
70c8708b
70cabd10
70880e12
700a704b
7b43bd10
7848b913
e0017809
78497808
2000ea41
7b434770
78c8b943
ea43788b
78482200
ea407809
e0072202
7808784a
78c9788b
2000ea42
2200ea43
2002ea41
00004770
4100f081
bf00e002
4300f083
ea4fb530
ea4f0441
ea940543
bf080f05
0f02ea90
ea54bf1f
ea550c00
ea7f0c02
ea7f5c64
f0005c65
ea4f80e2
ebd45454
bfb85555
dd0c426d
ea80442c
ea810202
ea820303
ea830000
ea800101
ea810202
2d360303
bd30bf88
4f00f011
3101ea4f
1c80f44f
3111ea4c
4240d002
0141eb61
4f00f013
3303ea4f
3313ea4c
4252d002
0343eb63
0f05ea94
80a7f000
0401f1a4
0e20f1d5
fa02db0d
fa22fc0e
1880f205
0100f141
f20efa03
fa431880
4159f305
f1a5e00e
f10e0520
2a010e20
fc0efa03
f04cbf28
fa430c02
18c0f305
71e3eb51
4500f001
f04fd507
f1dc0e00
eb7e0c00
eb6e0000
f5b10101
d31b1f80
1f00f5b1
0849d30c
0030ea5f
0c3cea4f
0401f104
5244ea4f
0f80f512
809af080
4f00f1bc
ea5fbf08
f1500c50
eb410000
ea415104
bd300105
0c4cea5f
eb414140
f4110101
f1a41f80
d1e90401
0f00f091
4601bf04
fab12000
bf08f381
f1a33320
f1b3030b
da0c0220
dd08320c
0c14f102
020cf1c2
f00cfa01
f102fa21
f102e00c
bfd80214
0c20f1c2
f102fa01
fc0cfa20
ea41bfdc
4090010c
bfa21ae4
5104eb01
bd304329
0404ea6f
da1c3c1f
dc0e340c
0414f104
0220f1c4
f004fa20
f302fa01
0003ea40
f304fa21
0103ea45
f1c4bd30
f1c4040c
fa200220
fa01f002
ea40f304
46290003
fa21bd30
4629f004
f094bd30
f4830f00
bf061380
1180f481
3d013401
ea7fe74e
bf185c64
5c65ea7f
ea94d029
bf080f05
0f02ea90
ea54d005
bf040c00
46104619
ea91bd30
bf1e0f03
20002100
ea5fbd30
d1055c54
41490040
f041bf28
bd304100
0480f514
f501bf3c
bd301180
4500f001
41fef045
0170f441
0000f04f
ea7fbd30
bf1a5c64
46104619
5c65ea7f
460bbf1c
ea504602
bf063401
3503ea52
0f03ea91
2100f441
bf00bd30
0f00f090
2100bf04
b5304770
6480f44f
0432f104
0500f04f
0100f04f
bf00e750
0f00f090
2100bf04
b5304770
6480f44f
0432f104
4500f010
4240bf48
0100f04f
bf00e73e
ea4f0042
ea4f01e2
ea4f0131
bf1f7002
437ff012
4f7ff093
5160f081
f0924770
bf140f00
4f7ff093
b5304770
7460f44f
4500f001
4100f021
bf00e720
0201ea50
4770bf08
f04fb530
e00a0500
0201ea50
4770bf08
f011b530
d5024500
eb614240
f44f0141
f1046480
ea5f0432
f43f5c91
f04faedc
ea5f0203
bf180cdc
ea5f3203
bf180cdc
eb023203
f1c202dc
fa000320
fa20fc03
fa01f002
ea40fe03
fa21000e
4414f102
bf00e6c1
f04fb570
f44c0cff
ea1c6ce0
bf1d5411
5513ea1c
0f0cea94
0f0cea95
f8def000
ea81442c
ea210603
ea23514c
ea50534c
bf183501
3503ea52
1180f441
1380f443
fba0d038
f04fce02
fbe10500
f006e502
fbe04200
f04fe503
fbe10600
f09c5603
bf180f00
0e01f04e
04fff1a4
7f00f5b6
7440f564
ea5fd204
416d0e4e
0606eb46
21c6ea42
5155ea41
20c5ea4f
505eea40
2eceea4f
0cfdf1b4
f5bcbf88
d81e6fe0
4f00f1be
ea5fbf08
f1500e50
eb410000
bd705104
4600f006
0101ea46
0002ea40
0103ea81
045cebb4
ebd4bfc2
ea41050c
bd705104
1180f441
0e00f04f
f3003c01
f11480ab
bfde0f36
f0012000
bd704100
0400f1c4
da353c20
dc1b340c
0414f104
0520f1c4
f305fa00
f004fa20
f205fa01
0002ea40
4200f001
4100f021
70d3eb10
f604fa21
0106eb42
0e43ea5e
ea20bf08
bd7070d3
040cf1c4
0520f1c4
f304fa00
f005fa20
f204fa01
0002ea40
4100f001
70d3eb10
0100f141
0e43ea5e
ea20bf08
bd7070d3
0520f1c4
f205fa00
0e02ea4e
f304fa20
f205fa01
0302ea43
f004fa21
4100f001
f204fa21
0002ea20
70d3eb00
0e43ea5e
ea20bf08
bd7070d3
0f00f094
f001d10f
00404600
0101eb41
1f80f411
3c01bf08
ea41d0f7
f0950106
bf180f00
f0034770
00524600
0303eb43
1f80f413
3d01bf08
ea43d0f7
47700306
0f0cea94
5513ea0c
ea95bf18
d00c0f0c
0641ea50
ea52bf18
d1d10643
0103ea81
4100f001
0000f04f
ea50bd70
bf060641
46194610
0643ea52
ea94d019
d1020f0c
3601ea50
ea95d113
d1050f0c
3603ea52
4610bf1c
d10a4619
0103ea81
4100f001
41fef041
0170f441
0000f04f
f041bd70
f44141fe
bd700178
f04fb570
f44c0cff
ea1c6ce0
bf1d5411
5513ea1c
0f0cea94
0f0cea95
f8a7f000
0405eba4
0e03ea81
3503ea52
3101ea4f
8088f000
3303ea4f
5580f04f
1313ea45
6312ea43
2202ea4f
1511ea45
6510ea45
2600ea4f
4100f00e
bf08429d
f1444296
f50404fd
d2027440
ea4f085b
1ab60232
0503eb65
ea4f085b
f44f0232
f44f1080
ebb62c00
eb750e02
bf220e03
46751ab6
000cea40
ea4f085b
ebb60232
eb750e02
bf220e03
46751ab6
005cea40
ea4f085b
ebb60232
eb750e02
bf220e03
46751ab6
009cea40
ea4f085b
ebb60232
eb750e02
bf220e03
46751ab6
00dcea40
0e06ea55
ea4fd018
ea451505
ea4f7516
ea4f1606
ea4303c3
ea4f7352
ea5f02c2
d1c01c1c
1f80f411
ea41d10b
f04f0100
f04f0000
e7b64c00
1f80f411
4301bf04
f1b42000
bf880cfd
6fe0f5bc
aeaff63f
0c03ebb5
ebb6bf04
ea5f0c02
f1500c50
eb410000
bd705104
4e00f00e
3111ea4e
045ceb14
ebd4bfc2
ea41050c
bd705104
1180f441
0e00f04f
e6903c01
0e06ea45
ea0ce68d
ea945513
bf080f0c
0f0cea95
af3bf43f
0f0cea94
ea50d10a
f47f3401
ea95af34
f47f0f0c
4610af25
e72c4619
0f0cea95
ea52d106
f43f3503
4610aefd
e7224619
0641ea50
ea52bf18
f47f0643
ea50aec5
f47f0441
ea52af0d
f47f0543
e712aeeb
d211004a
1200f512
d50dd211
7378f46f
5262ebb3
ea4fd40e
f04323c1
ea434300
fa235350
4770f002
0000f04f
ea504770
d1023001
30fff04f
f04f4770
47700000
4000f080
bf00e002
4100f081
bf1f0042
0341ea5f
0f03ea92
6c22ea7f
6c23ea7f
ea4fd06a
ebd26212
bfc16313
404118d2
40414048
425bbfb8
bf882b19
f0104770
f4404f00
f0200000
bf18407f
f0114240
f4414f00
f0210100
bf18417f
ea924249
d03f0f03
0201f1a2
fc03fa41
000ceb10
0320f1c3
f103fa01
4300f000
4249d502
0040eb60
0f00f5b0
f1b0d313
d3067f80
ea4f0840
f1020131
2afe0201
f1b1d251
eb404f00
bf0850c2
0001f020
0003ea40
00494770
0000eb40
0f00f410
0201f1a2
fab0d1ed
f1acfc80
ebb20c08
fa00020c
bfaaf00c
50c2eb00
43184252
40d0bfbc
47704318
0f00f092
0100f481
f480bf06
32010000
e7b53b01
0341ea4f
6c22ea7f
ea7fbf18
d0216c23
0f03ea92
f092d004
bf080f00
47704608
0f01ea90
2000bf1c
f0124770
d1044f7f
bf280040
4000f040
f1124770
bf3c7200
0000f500
f0004770
f0434300
f44040fe
47700000
6222ea7f
4608bf16
6323ea7f
02424601
ea5fbf06
ea902341
f4400f01
47700080
0300f04f
bf00e004
4300f010
4240bf48
0c00ea5f
4770bf08
4396f043
f04f4601
e01c0000
0201ea50
4770bf08
0300f04f
bf00e00a
0201ea50
4770bf08
4300f011
4240d502
0141eb61
0c01ea5f
4684bf02
20004601
43b6f043
f1a3bf08
f5a35380
fabc0300
3a08f28c
53c2eba3
fa01db10
4463fc02
fc02fa00
0220f1c2
4f00f1bc
f202fa20
0002eb43
f020bf08
47700001
0220f102
fc02fa01
0220f1c2
004cea50
f202fa21
0002eb43
ea20bf08
477070dc
0cfff04f
52d0ea1c
ea1cbf1e
ea9253d1
ea930f0c
d06f0f0c
ea80441a
02400c01
ea5fbf18
d01e2141
6300f04f
1050ea43
1151ea43
3101fba0
4000f00c
0f00f5b1
0049bf3e
71d3ea41
ea40005b
f1620001
2afd027f
f1b3d81d
eb404f00
bf0850c2
0001f020
f0904770
f00c0f00
bf084c00
ea4c0249
ea402050
3a7f2051
f1d2bfc2
ea4003ff
477050c2
0000f440
0300f04f
dc5d3a01
0f19f112
f000bfdc
47704000
0200f1c2
fa210041
f1c2f102
fa000220
ea5ffc02
f1400031
ea530000
bf08034c
70dcea20
f0924770
f0000f00
bf024c00
f4100040
3a010f00
ea40d0f9
f093000c
f0010f00
bf024c00
f4110049
3b010f00
ea41d0f9
e78f010c
53d1ea0c
0f0cea92
ea93bf18
d00a0f0c
4c00f030
f031bf18
d1d84c00
0001ea80
4000f000
f0904770
bf170f00
4f00f090
f0914608
f0910f00
d0144f00
0f0cea92
0242d101
ea93d10f
d1030f0c
bf18024b
d1084608
0001ea80
4000f000
40fef040
0000f440
f0404770
f44040fe
47700040
0cfff04f
52d0ea1c
ea1cbf1e
ea9253d1
ea930f0c
d0690f0c
0203eba2
0c01ea80
ea4f0249
d0372040
5380f04f
1111ea43
1310ea43
4000f00c
bf38428b
f142005b
f44f027d
428b0c00
1a5bbf24
000cea40
0f51ebb3
eba3bf24
ea400351
ebb3005c
bf240f91
0391eba3
009cea40
0fd1ebb3
eba3bf24
ea4003d1
011b00dc
ea5fbf18
d1e01c1c
f63f2afd
428baf50
50c2eb40
f020bf08
47700001
4c00f00c
2050ea4c
bfc2327f
03fff1d2
50c2ea40
f4404770
f04f0000
3a010300
f092e737
f0000f00
bf024c00
f4100040
3a010f00
ea40d0f9
f093000c
f0010f00
bf024c00
f4110049
3b010f00
ea41d0f9
e795010c
53d1ea0c
0f0cea92
0242d108
af7df47f
0f0cea93
af70f47f
e7764608
0f0cea93
024bd104
af4cf43f
e76e4608
4c00f030
f031bf18
d1ca4c00
4200f030
af5cf47f
4300f031
af3cf47f
bf00e75f
3cfff04f
bf00e006
0c01f04f
bf00e002
0c01f04f
cd04f84d
0240ea4f
0341ea4f
6c22ea7f
ea7fbf18
d0116c23
ea52b001
bf180c53
0f01ea90
ebb2bf58
bf880003
bf3817c8
70e1ea6f
f040bf18
47700001
6c22ea7f
ea5fd102
d1052c40
6c23ea7f
ea5fd1e4
d0e12c41
0b04f85d
bf004770
46084684
e7ff4661
f7ffb50f
2800ffc9
f110bf48
bd0f0f00
ed08f84d
fff4f7ff
2001bf0c
f85d2000
bf00fb08
ed08f84d
ffeaf7ff
2001bf34
f85d2000
bf00fb08
ed08f84d
ffe0f7ff
2001bf94
f85d2000
bf00fb08
ed08f84d
ffd2f7ff
2001bf94
f85d2000
bf00fb08
ed08f84d
ffc8f7ff
2001bf34
f85d2000
bf00fb08
0240ea4f
4ffef1b2
f04fd30f
ebb3039e
d90d6212
2300ea4f
4300f043
4f00f010
f002fa23
4240bf18
f04f4770
47700000
0f61f112
0242d101
f010d105
bf084000
4000f06f
f04f4770
47700000
d20e0042
4ffef1b2
f04fd30b
ebb3039e
d4096212
2300ea4f
4300f043
f002fa23
f04f4770
47700000
0f61f112
0242d101
f04fd102
477030ff
0000f04f
bf004770
e92d2a0f
f24003f0
ea418095
079b0300
8092f040
6004680c
6045684d
f1a2688e
60860310
461d68cc
60c42d0f
1600f3c3
0410f101
0310f100
b166d922
601e6826
605e6866
609e68a6
3d1068e6
341060de
2d0f3310
6826d914
6866601e
68a6605e
68e6609e
692660de
6966611e
69a6615e
69e6619e
61de3d20
33203420
d8ea2d0f
0310f1a2
040ff023
030ff002
2b033410
0804eb00
d9514421
0904f1a3
ea4f460b
eb010999
f8530c89
ebc16b04
4644050c
0c04f10c
f8444563
f3c56b04
d0120580
f853b12d
45635b04
5b04f844
461ed00b
f8564625
f8457b04
685f7b04
60671d33
45631d2c
f109d1f3
009c0301
f0021909
44440203
4623b1da
f803780d
18a25b01
191443e4
f0044293
d0100401
f811b12c
f8034f01
42934b01
784dd009
f804461c
788d5b01
1c63705d
42933102
e8bdd1f5
477003f0
e7dd4604
e7dc4604
461a4644
bf00e7d8
0784b4f0
f0004603
1e54808e
f0002a00
07e58088
d411b2ce
1e67461a
6b01f802
46154613
d00f0792
d07a2c00
6b01f803
463c079a
d007461d
e7ed3c01
f8034603
079a6b01
d1f7461d
d9522c03
ea46b2ce
2c0f2706
4307ea47
f1a4d92d
46170210
f3c22f0f
602b1600
60ab606b
f10560eb
d9160210
3f10b13e
60536013
60d36093
2f0f3210
3f20d90d
0610f102
60536013
60d36093
61536113
61d36193
2f0f3220
f1a4d8f1
f0220210
f004020f
3210040f
44152c03
1f27d91d
462a463e
f8422e03
f3c73b04
d90d0780
3e04b127
f8422e03
d9073b04
3e084617
3b04f847
1d3a6053
d8f72e03
f0231f23
1d130203
0403f004
b1b418ed
b2c9462b
1b01f803
43ed192c
42a31962
0501f002
b11dd00b
1b01f803
d00642a3
f802461a
70591b01
42a31c53
bcf0d1f8
46054770
e78d4614
00000000
3441f19a
4a003d52
