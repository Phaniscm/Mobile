0004909c
544f4f42
52455620
382e3020
0000332e
00000000
00000000
00000000
0804909c
00040404
00040404
0804ae9c
00040404
00040404
00040404
00040404
00040013
00040013
0804ba9c
00040013
0804b69c
00040013
00040013
00040013
0804989c
00040404
00040404
0804909c
00040404
00040404
00040404
00040404
0804909c
0804959c
00040404
00040404
00040404
00040404
00040404
00040404
fff30004
00040404
00040404
00040404
00040404
00040404
00040404
00040404
00040013
00040013
00040404
00040404
00040404
00040404
00040404
00040404
fff30004
00040404
00040404
00040404
00040404
00040404
00040404
00040404
00040013
00040013
00040404
00040404
00040404
00040404
00040404
00040404
0001c800
0001d5e8
00000000
04081000
66001100
000000ff
0f0e270c
1817160a
08070625
0e0d0c09
230b0a0f
07062524
37360908
35343938
0633302f
25090807
15292827
11181716
39383736
0a0a0909
09090909
09090904
0a0a0909
0909090a
09090409
04040909
09090404
09090909
09090909
09090909
09090909
09090909
0504ff03
ffffff02
01010109
04040301
09020205
01010909
0d0d0101
0d0d0e0e
010c0b0b
09010101
ffffffff
05ffffff
0e0e0d0d
0011cafc
0011cb00
0011cb2c
0011cba4
0011cbb0
0011cbb8
0011cbc0
0011cbdc
0011cbfc
001179e4
00117a6c
00117aa4
001179bc
001187a8
00117cb0
0010c4fc
0010c1bc
0010c1c8
0010c1cc
0010c1fc
0010c20c
001187f8
0010c684
0010c1b8
0010c1f8
0010c1c0
0010c1c4
0010c278
00180004
00180004
000014ac
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
0580301c
4130311c
60076c0c
60060815
4140311c
211c4006
4c0f0040
311c6286
6c0c4105
0140341c
0140331c
60060394
f01c3464
f11cbc00
0ebc0001
00130850
00000804
00000004
08040013
08040013
b400f01c
0001f11c
080746bc
00000804
7f36ff16
082868bc
ff56fe76
ff160404
68bc7f36
fe760828
0404ff56
7f36ff16
0807cabc
ff56fe76
00130404
00130464
00000804
8624301c
2404311c
251c4c0c
4c0f0018
301c6c0c
311c0094
6c0c4080
0014033c
00000804
211c4006
62060001
4600311c
303c4c0f
2086200c
4613111c
0c0b6c80
311c6286
4c0f4600
08040364
600620c3
4140311c
011c0006
0c0f0200
111c2006
68802010
080c133c
640e6006
011c0006
6800104e
100c233c
6472680c
640b680f
65723364
0004640e
003c040b
08040b4b
0136f016
60c3fe96
42c381c3
0240503c
323c412c
67d21004
1a4b323c
305c3264
03336ee7
17548007
0580101c
4130111c
740f640c
6872612c
08c3612f
24d1705c
241c27c3
323c0007
792f1a5b
6ee7265c
640f740c
303c192c
60071004
365c2a54
60276ee4
301c0994
311c800c
4c0c4600
0700251c
604703b3
301c0994
311c800c
4c0c4600
0600251c
7f850273
0ab46027
800c201c
4600211c
351c680c
680f5000
301c0113
311c800c
4c0c4600
4c0f4a72
6e04165c
1004313c
301c69f2
311cc800
4c0c0001
800742a3
365c3254
22866ee4
4105111c
0804203c
1b946007
53c3640c
301c5364
311cc828
6c0c0001
245c48c3
145c2473
745c2483
e0370784
0761045c
435c0077
02c314e4
32c34026
01934664
53c3640c
353c5364
7bd20384
353c45d2
608718cb
565cf654
18b36e07
32c3596c
4001701c
1000711c
47c33783
095434e4
0014313c
16946007
0014323c
12546007
c828301c
0001311c
335c6c0c
06c321a4
366418c3
8048201c
4600211c
6072680c
192c680f
1004303c
3b546007
1a4b703c
6ee7765c
111c2286
e0074105
08c32294
0564305c
1004533c
c828201c
0001211c
680caed2
0784105c
205c2037
40770764
06c38c4c
27c318c3
013337c3
a037680c
8c4ca077
18c306c3
35c325c3
0e734664
23c3640c
323c2364
7bd20384
0121365c
60076732
323c6854
608718cb
0c73f254
375c78c3
133c0564
201c1004
211cc828
2ad20001
303c480c
075c09cb
00370784
0764175c
480c00b3
09cb303c
20772037
06c3884c
402618c3
62864664
4105311c
33646c0c
6e07365c
0121265c
63324732
341c44d2
01730003
236423c3
0074323c
6ee7365c
05356067
0044323c
6ee7365c
6ee4365c
0e946087
c828301c
0001311c
335c6c0c
03c60484
04f23664
065c00a6
265c6ee7
792c6ee4
1a5b323c
792f6872
22e6101c
4c097880
540c48f2
0580301c
4130311c
00f34c0f
0580301c
4130311c
740f6c0c
80760296
08040f56
24b1315c
13946b47
cf30301c
0001311c
4e4d4b26
c828301c
0001311c
335c6c0c
015c0424
115c24b9
366424c3
00000804
40c31016
6e29205c
341c32c3
60070001
620c1c54
205c7112
6d002764
f000321c
331c6c0b
11945aa5
cf30301c
0001311c
4f6d4b26
c828301c
0001311c
335c6c0c
103c0a04
36640340
6e29245c
341c32c3
60070002
345c1e54
71122ba4
5104245c
321c6d00
6c0bf000
5aa5331c
301c1294
311ccf30
4b260001
301c4f8d
311cc828
6c0c0001
0a04335c
143c04c3
36645680
08040856
0136f016
70c3ff96
200761c3
80c35954
0df8821c
c828501c
0001511c
315c540c
001c25c4
2c00f000
7112786c
15a4425c
258008c3
46644706
365c540c
001c25c4
2c00f400
7112786c
15a4425c
8000001c
0001011c
201c2580
46640c00
175c740c
203771a4
0e64435c
268608c3
32c34006
30c34664
275c8006
02c37164
169430e4
6e6c740c
16c307c3
40c33664
2222031c
031c0454
0a945555
c828301c
0001311c
6e8c6c0c
16c307c3
301c3664
311cc828
6c0c0001
07c36dec
24c316c3
01963664
0f568076
00000804
a5063016
4110511c
c828401c
0001411c
341c740b
7dd20002
6d8c700c
ff333664
08040c56
313c200c
66d20014
6186404c
4140311c
313c4c0f
66d20044
6286408c
4140311c
313c4c0f
66d20084
6a0640ac
4140311c
08044c0f
313c1016
60070024
301c3f54
311c0480
4c0c4130
4c0f4172
211c4686
680c4140
0040341c
40c97dd2
40e942c3
422c323c
8028201c
4113211c
313c680e
60070014
60891c54
60a943c3
422c233c
8024301c
4113311c
81094c0e
812914c3
40ac243c
4c0e6105
31c32149
213c2169
301c41ac
311c8030
4c0e4113
211c4686
680c4140
0040341c
08567dd2
00000804
fe961016
c828401c
0001411c
4037900c
445c6077
402614e4
466432c3
08560296
00000804
08d43cbc
00000804
001c3016
011cd800
405c0001
8bd26e29
0014343c
d834501c
0001511c
521c6ff2
01930534
c828301c
0001311c
6f2c6c0c
201c14c3
366400fa
301c54c3
311c0580
6c0c4130
111c2006
31831000
301c6ed2
311ccf30
4b260001
0115235c
c800301c
0001311c
2c0f2026
c800401c
0001411c
6007700c
301c2194
311cc828
6c0c0001
0444335c
00073664
255c1754
40272469
301c1394
311cd800
335c0001
341c6e04
6ad20001
cf30301c
0001311c
135c2b26
500f011d
40060053
c828301c
0001311c
335c6c0c
001c2044
011cd800
15c30001
301c3664
311cc800
4c0c0001
35944007
d800101c
0001111c
6e04315c
0100341c
2b946007
cf30301c
0001311c
235c4b26
315c0125
60476ee4
60870554
60270354
301c0e94
311cc828
6c0c0001
07a4335c
d800001c
0001011c
0e533664
035460a7
6e946007
c828301c
0001311c
335c6c0c
000607e4
0c933664
2441355c
262664f2
2445155c
45544007
d800001c
0001011c
31c3216c
4001341c
4001331c
301c3a94
311ccf30
4b260001
012d235c
311c6006
13831000
12542007
c828301c
0001311c
335c6c0c
15c321a4
201c3664
211c8048
680c4600
680f6072
255c0173
323c2449
758002c7
0f84235c
04bc43d2
301c0843
311cc828
6c0c0001
2449255c
001c8fac
011cd800
155c0001
60062441
03134664
cf30301c
0001311c
135c2b26
301c0135
311cc828
6c0c0001
2449255c
001c8fac
011cd800
155c0001
60062441
00134664
08040c56
13640364
0104303c
68d22312
311c60c6
45804080
ffef041c
604600b3
4080311c
60264580
33643023
0804680e
313c1364
4486080c
4080211c
640b2d00
40263364
000d023c
328320e3
0804640e
111c2f86
40064010
4010211c
341c640b
63d20008
ff73680b
00000804
8157f016
71c30364
52c37364
63c35364
89f26364
311c6206
20264020
60452c0e
06532c0e
0ff4343c
211c4006
6d002010
080c233c
00c13f5c
343c680e
2006420b
2010111c
233c6c80
2197080c
420b313c
343c680e
6007808c
341c1754
400600ff
2010211c
233c6d00
313c080c
680e440b
c08c343c
211c4006
6d002010
080c233c
783231c3
2186680e
4010111c
0080301c
4006640e
6206440e
4010311c
61064c0e
4010311c
4c0e4826
ac0e6f05
cc0e6085
0080301c
203c640e
60060ff4
4010311c
203c4c0e
6085408c
321c4c0e
ec0e00bc
a40ea006
440e4066
08040f56
301cfe96
311cd800
335c0001
60076ee4
4f861594
4010211c
3364680b
00363f5c
00333f5c
0008341c
600678d2
4010311c
23c36c0b
40372264
301c0173
0c0c0b00
0200101c
08c65ebc
326430c3
3f5c6037
03c30001
08040296
30c3fe96
60373264
d800301c
0001311c
6ee4335c
13946007
311c6006
40174010
42864c0e
4010211c
3364680b
00363f5c
00333f5c
0040341c
00d378d2
00013f5c
0abc03c3
02960861
00000804
50c3f016
63c342c3
0c064006
41e4e066
6c861b14
1530141d
141d0412
33643100
233c780e
313cc187
141d3e87
69803300
23c36612
301c2364
141d03e8
41573230
0006680e
40470233
313c0994
141d080c
303c1370
0180088c
21320073
40250112
d6944147
0f561fe6
00000804
600620c3
4140311c
011c0006
0c0f0200
111c2006
68802010
080c133c
640e6006
011c0006
6800104e
100c233c
6472680c
640b680f
351c3364
640e0420
3364640b
00c0351c
0804640e
211c4006
6100104e
100c233c
6492680c
4006680f
2010211c
61126100
4c0e4406
00000804
3f36f016
d0c3fd96
a2c3c1c3
93c3a364
40069364
00562f5c
00462f5c
60776006
0397a106
12540007
51c32397
00ff541c
0454a107
26bc0106
0397080a
420b303c
04546127
26bc0126
2ac3080a
12544007
211c4286
680c4105
0038341c
931c6bd2
a4dc0001
680c0011
18cb333c
44dc6087
401c0011
411cc828
700c0001
05c36c2c
20063664
2010111c
733c7480
b01c080c
b11c0014
801c4105
811c0000
2ac34040
10544007
600c0bc3
0038341c
931c6bd2
24dc0001
600c000f
18cb333c
c4dc6087
001c000e
011cffff
38c3000f
7c0c0c0f
7c0f6b72
640c1bc3
0ac35c0c
14540007
0038341c
10546007
0001931c
0bc30794
333c600c
608718cb
60060754
4040311c
4c2f4806
32c31933
1000341c
e3546007
38c30026
7c0c0c2f
7c0f6b72
2bc32046
5c0c680c
00070ac3
341c1454
60070038
931c1054
07940001
600c0bc3
18cb333c
07546087
311c6006
28064040
14932c2f
341c32c3
60071000
7c0ce354
2000341c
0014213c
189432e4
00534006
18c34026
6077640c
001c6057
011cffff
61a0000f
60576077
f49430e4
640f18c3
642f6026
ed544007
7c0cf2f3
7c0f6b72
20a72025
4806bf94
442f18c3
6077640c
001c6057
011cffff
61a0000f
40066077
323c0193
23c30010
101c2364
111cffff
31c30000
055423e4
341c7c0c
72d21000
fff0323c
001c3364
011cfffd
10c30000
a9dc31e4
c057fff6
c828301c
0001311c
0dc34c0c
6ea4105c
6ec4405c
00803f3c
a80c6037
14c301c3
3f3c26c3
566400a0
00531f5c
325c2cc3
31e42473
2f5c0894
0cc30043
2483305c
0c5423e4
c828201c
0001211c
8eec680c
2f5c0dc3
3cc30043
001c4664
011cc828
600c0001
0a84435c
00530f5c
00431f5c
63d74397
101c4664
111cc828
640c0001
1504335c
36640aa6
c828201c
0001211c
035c680c
06641524
326430c3
64dc6aa7
0396fff0
0f56fc76
00000804
311c6006
40264140
301c4c0f
311c4240
141d000f
23c33030
301c2364
311c0084
4c0e4040
60852006
301c2c0e
141d03e8
23c33030
301c2364
311c008c
4c0e4040
2c0e6085
00000804
0f36f016
80c3fd96
63c371c3
0184af5c
c828401c
0001411c
335c700c
0ac315a4
420612c3
b01c3664
b11cfab8
94c30001
631c56c3
03351000
1000501c
3bc3daa0
19c34c0c
335c640c
023c0904
208601c0
ea58201c
0001211c
29c33664
a037680c
20772026
8cec20b7
17c308c3
8000201c
0001211c
ea58301c
0001311c
3bc34664
19c34c0c
335c640c
023c0904
214601c0
e640201c
0001211c
29c33664
af5c680c
8ccc0007
8000001c
0001011c
201c1ac3
211ce640
35c30001
fe804664
c0078584
0396b894
0f56f076
00000804
fd96f016
71c360c3
13c352c3
30c3082b
0020361c
7f327fe5
080c033c
542900b7
0014323c
323c66f2
63f20044
00b70272
c828301c
0001311c
20376c0c
40774217
16e4435c
00413f5c
16c303c3
353c27c3
46640080
0f560396
00000804
fa967016
42c350c3
4c2b03c3
361c32c3
7fe50020
233c7f32
4177080c
63d26317
41774472
323c4029
67f20014
0044323c
c15764f2
c177c272
c828301c
0001311c
303c4c0c
60370080
60776297
601c80b7
611cfacc
c0f70001
613762d7
1704425c
00a16f5c
25c306c3
46646006
0e560696
00000804
1f36f016
80c3fd96
93c371c3
cf5cc357
af5c01c4
401c01e4
411cc828
700c0001
15a4335c
12c30cc3
36644206
56c3b4c3
1000631c
501c0335
daa01000
69d23ac3
680c2bc3
af5ca037
40260027
011340b7
680c2bc3
af5ca037
af5c0027
8cec0047
17c308c3
8000201c
0001211c
466439c3
680c2bc3
0007cf5c
001c8ccc
011c8000
1cc30001
35c329c3
c4d24664
8584fe80
0396f9f3
0f56f876
00000804
fc967016
c21743c3
ce58501c
0001511c
6bd27409
61e74006
133c0654
20f70010
00612f5c
0773540d
041c01c3
0af2f000
6e0068a0
ffff401c
0000411c
32e424c3
301c17b4
311cc828
6c0c0001
21e4335c
25a4265c
80262037
20068077
8e0c20b7
13c302c3
1ac0263c
46646406
301c0313
311cc828
6c0c0001
21e4335c
25a4265c
80262037
00b78077
02c38e0c
263c13c3
301c1ac0
466400d8
340d2026
0e560496
00000804
40c37016
201c61c3
211cbaad
205c0000
301c6f87
311cc828
6c0c0001
15a4535c
c830301c
0001311c
6f64205c
145c0d00
26c36f44
345c5664
6f006f64
6f67345c
900d301c
0000311c
6f87345c
08040e56
1f36f016
50c3fc96
b2c361c3
705cc3c3
301c6fa4
311cce54
6c0c0001
600760f7
001584dc
ce4c301c
0001311c
ce0c101c
0001111c
301c2c0f
311cc828
6c0c0001
15a4335c
155c01c3
48066f44
2f5c3664
32c30061
0294c847
a3c36026
363ca264
333c0346
7fe50b0d
f88c833c
98a39ac3
6df239c3
0b54c567
0954c4a7
0754ca27
0554c4c7
c54719c3
001294dc
341c744c
60071000
000aa2dc
c828301c
0001311c
335c6c0c
101c1584
14800df8
36642706
0564375c
211c4006
32830200
23546007
0554ca27
0354c4c7
0f94c547
0c04375c
f000401c
301c4e00
311cce4c
6c0c0001
68a02c2c
04933483
0c04375c
efc0101c
301c4c80
311cce0c
8c4c0001
28056a20
05d33183
0554ca27
0354c4c7
1a94c547
233c7c6c
301c880c
311cce4c
6c0c0001
68a02c2c
c000321c
f000201c
355c3283
301c7027
311cce0c
80060001
8c4f8c8f
7c6c0233
880c233c
ce0c301c
0001311c
68a02c4c
bfc0321c
f000201c
355c3283
401c7027
411cce0c
704c0001
7047355c
155c308c
500b7067
6ff6255c
355c706c
314c7127
7147155c
c828301c
0001311c
335c6c0c
201c15a4
15000e14
0180143c
36644206
355c70ac
055c7087
48c37024
8ef22046
60262ac3
10944007
c5672206
64060754
0a54c4a7
0594ca27
155c2106
02136fe6
0594c4c7
355c6126
01536fe6
c5472146
fe930794
ce0c301c
0001311c
363c0c8c
333c0256
7fe50b0d
f88c233c
62f238c3
744c45d2
0c4b333c
744c0093
0bcb333c
4b546007
02b6363c
0b0d333c
133c7fe5
46f2f88c
49c325f2
15948007
400707d3
375c1254
101c2824
111cbbbb
21c30000
339432e4
ce0c301c
0001311c
475c6c6c
04b32944
18542007
26a4375c
aaaa401c
0000411c
31e414c3
301c2094
311cce0c
6c6c0001
27c4275c
34e442c3
20261634
7187155c
3c3c0253
7d8002c7
1e80233c
ce0c301c
0001311c
880c6c6c
31e414c3
40260434
7187255c
ce0c201c
0001211c
888c684c
7c6c4e00
74126332
23e47fe5
40260435
7187255c
00d310c3
6f64305c
6f24405c
b55c2e00
155c6f67
355c6f27
68d27184
900d101c
0000111c
6f87155c
201c05d3
211cbaad
255c0000
301c6f87
311cce54
0c0c0001
1c940007
fff4313c
18546007
c828301c
0001311c
335c6c0c
275c21e4
401c25a4
1483f000
20262037
00b72077
02c38e0c
273c13c3
64061ac0
64064664
4110311c
4c0e4046
ce54301c
0001311c
40254c0c
04964c0f
0f56f876
00000804
40c33016
60cc51c3
211c4006
32830010
305c6ed2
7fe56ee4
09b46027
c828301c
0001311c
335c6c0c
36640804
6fa7545c
9000301c
0001311c
6f47345c
900d201c
0000211c
6f87245c
345c6006
0c566f67
00000804
3f36f016
81c3fe96
c3c3d2c3
20c30449
903c0469
0006412c
01a11f5c
361c31c3
7fe50002
b33c7f32
201ca80c
211cc828
680c0001
15a4335c
303c6037
48c3180c
233c7180
2c29061e
412c213c
243c8c49
2c69812c
c12c213c
3cc349c3
25c4335c
703c3180
373c0010
48c3180c
56c3d180
009e353c
7c9d043c
402c433c
46c38077
0d003bc3
28802dc3
a3c36057
011e343c
852c233c
36646017
103c08c3
14097c9d
40ac303c
213c3009
786981ac
64f26732
07c39284
0296f773
0f56fc76
00000804
3f36f016
50c3f396
c2c391c3
6f5c60f7
001c0301
14001258
44490137
446932c3
41acb23c
c828401c
0001411c
335c700c
0f3c15a4
201c0140
350022bc
36644206
0000a01c
0026363c
7f327fe5
a80cd33c
00101a3c
180c313c
518049c3
1c9d043c
082940c3
422c303c
613c2849
801c81ac
3a3c0000
29c3180c
733c6980
56c300c0
1000631c
501c03f4
daa01000
c828401c
0001411c
1bc3700c
005c00d7
440025c4
2026a037
20b72077
3cc38cec
0b840cc3
201c2d00
211c8000
61170001
401c4664
411cc828
700c0001
15a4435c
10c31c09
303c1c29
3c4940ac
81ac313c
323c5c69
08c3c1ac
1dc36180
101c0c80
111c8000
25c30001
b5844664
03f4c007
f8138584
00101a3c
180c313c
718049c3
67326c69
a1c363f2
0d96f3d3
0f56fc76
00000804
0336f016
fbd0f21c
31c380c3
921c90c3
29c322b8
331c080c
14dc2222
301c000b
311cce50
6c0c0001
92dc6007
703c000a
341c01c0
60070001
401c3054
411cc828
700c0001
08e4335c
202607c3
20c33664
6f3c700c
335c0080
06c315a4
201c12c3
36640428
2f5c4106
700c0045
08e4335c
210607c3
50c33664
19c3700c
101c440c
20370428
5aa5101c
435c2077
08c30964
25c312c3
466436c3
ce50301c
0001311c
341c6c0c
60070002
401c3254
411cc828
700c0001
08e4335c
204607c3
20c33664
6f3c700c
335c0080
06c315a4
201c12c3
36640428
2f5c4126
700c0045
08e4335c
212607c3
50c33664
38c3500c
22b8321c
101c6c0c
20370428
5aa5101c
425c2077
08c30964
25c313c3
466436c3
ce50301c
0001311c
341c6c0c
60070004
401c3054
411cc828
700c0001
08e4335c
206607c3
20c33664
6f3c700c
335c0080
06c315a4
470612c3
41463664
00452f5c
335c700c
07c308e4
36642146
500c50c3
321c38c3
6c0c22b8
20372706
5aa5101c
425c2077
08c30964
25c313c3
466436c3
ce50301c
0001311c
4c0f4006
0430f21c
0f56c076
00000804
0136f016
80c3f896
52c371c3
c828601c
0001611c
401c780c
411c9000
335c0001
04c31584
0400101c
b00f3664
ce50301c
0001311c
6ad26c0c
2222531c
780c0794
04a4335c
15c308c3
501c3664
511cc828
740c0001
21e4235c
1ac0673c
25a4175c
71127c6c
f000321c
60266037
60066077
8a0c60b7
12c301c3
640626c3
740c4664
21e4235c
25a4175c
71127c6c
f000321c
301c6037
311c9000
60770001
0400301c
301c60b7
3f5c0100
60060066
60266137
60066177
61f761b7
01c38a2c
26c312c3
46646046
235c740c
175c21e4
7c6c25a4
321c7112
6037f400
8000301c
0001311c
301c6077
60b70c00
0100301c
00663f5c
61376006
61776026
61b76006
8a2c61f7
12c301c3
604626c3
08964664
0f568076
00000804
0f36f016
40c3f896
a0c351c3
0df8a21c
c828701c
0001711c
205c7c0c
403771a4
0e64635c
26860ac3
32c34006
045c6664
b01c7167
b11c8000
5c0c0001
25c4355c
f400001c
746c2c00
425c7112
0bc315a4
201c2580
46640c00
235c7c0c
953c21e4
155c1ac0
746c25a4
321c7112
6037f000
0001801c
00278f5c
80b78006
01c3ca0c
29c312c3
66646406
235c7c0c
155c21e4
746c25a4
321c7112
6037f000
0027af5c
60b76706
0100a01c
0066af5c
8f5c8137
81b700a7
ca2c81f7
12c301c3
604629c3
7c0c6664
21e4235c
25a4155c
7112746c
f400321c
bf5c6037
001c0027
00b70c00
0066af5c
8f5c8137
81b700a7
8a2c81f7
12c301c3
604629c3
08964664
0f56f076
00000804
0336f016
fcf8f21c
61c372c3
23c36264
323c2264
833cfff0
18c3f88c
231c28f2
055400f1
00f2231c
000fc4dc
1c80973c
c828501c
0001511c
105c740c
203771a4
0e64435c
101c09c3
400602e4
466432c3
2567075c
25c4175c
1154c007
121c540c
7c6cf400
425c7112
001c15a4
011c8000
25800001
0c00201c
02134664
475c740c
460025e4
15a4335c
8000001c
0001011c
4000123c
0c00201c
08c33664
6a540007
02008f3c
c828501c
0001511c
275c740c
335c25e4
08c315a4
25c4475c
201c2a00
366402e8
235c740c
673c21e4
175c1ac0
7c6c25a4
321c7112
6037e000
00770026
60b76006
01c38a0c
26c312c3
46646406
235c740c
175c21e4
7c6c25a4
321c7112
6037e000
00278f5c
02e8401c
001c80b7
0f5c0100
60060066
80266137
61b78177
8a2c61f7
12c301c3
604626c3
740c4664
21e4235c
25a4175c
71127c6c
e400321c
001c6037
011c8000
00770001
0c00301c
401c60b7
4f5c0100
00060066
60260137
01b76177
8a2c01f7
12c301c3
604626c3
501c4664
511cc828
740c0001
21e4235c
1ac0673c
25a4375c
25e4475c
00268037
20060077
8a0c20b7
12c303c3
640626c3
740c4664
21e4335c
25a4275c
25e4475c
9f5c8037
001c0027
00b702e8
0100101c
00661f5c
81378006
01770026
81f781b7
02c38e2c
26c313c3
46646046
235c740c
175c21e4
375c25a4
321c25e4
60370400
8000301c
0001311c
401c6077
80b70c00
0100001c
00660f5c
61376006
81778026
61f761b7
01c38a2c
26c312c3
46646046
0308f21c
0f56c076
00000804
3f36f016
70c3ee96
205c21b7
40876fe3
301c1e94
311cc828
6c0c0001
71a4175c
435c2037
001c0e64
011c8000
101c0001
40060c00
466432c3
5555201c
7084475c
05e454c3
004504dc
00045b9c
d21cd7c3
323c0e40
7fe50106
f88c633c
fff0323c
60273364
c4f20535
24dc4407
61970021
25c4935c
7024875c
7044a75c
0206323c
033c7fe5
323cf88c
7fe50026
f88c133c
7c4c10a3
233c29d2
533c0c4b
7c8c0c8b
0b0b433c
233c00f3
533c0bcb
433c0c0b
40070b8b
61971a54
221c23c3
0ef20508
20c30197
04d8221c
375cc9f2
333c7004
321c02c7
c19701c8
375c5980
090c7124
36e460c3
004000dc
375c0ac3
41807064
786cc197
74126832
23e47fe5
003f45dc
275ca9d2
32c36ff3
0008341c
b2dc6007
89d2003e
6ff3475c
341c34c3
60070004
003e22dc
6ff3575c
041c05c3
04f20008
b0c30237
401c0cd3
411cc828
601c0001
bf0022b8
2d542007
b21cb7c3
700c1ea0
335c540c
023c0904
212601c0
36642bc3
1ea4101c
375cdc80
580c7144
30e402c3
700c4435
335c540c
023c0904
204601c0
36642bc3
7144375c
21c3380c
b4dc32e4
301c003a
311cce50
4c0c0001
05934172
b21cb7c3
700c1a88
335c540c
023c0904
210601c0
36642bc3
1a8c001c
375cdc00
380c7144
32e421c3
700c1835
335c540c
023c0904
202601c0
36642bc3
7144375c
54c3980c
f4dc35e4
301c0037
311cce50
4c0c0001
4c0f4072
d8cb6bc3
a6a4c237
18c38984
c83c98c3
601c0400
611cce0c
501c0001
511cc828
740c0001
15a4335c
480606c3
275c3664
32c36ff3
0004341c
92dc6007
540c000a
22b8401c
6c0c7e00
0904425c
01c0033c
2dc32146
740c4664
1584335c
0180063c
36642206
03808f3c
22bc001c
03771c00
335c740c
08c315a4
42062357
740c3664
00078f5c
06c38ccc
2dc318c3
46646806
6ff3175c
341c31c3
6fd20002
af5c740c
8f5c0007
40060027
8cac40b7
1cc302c3
3dc328c3
01534664
8f5c740c
8ccc0007
18c30cc3
3ac32dc3
493c4664
81f70180
c828601c
0001611c
335c780c
08c315c4
420614c3
00073664
580c6454
22b8501c
6c0c7e80
0904425c
01c0033c
2dc32066
780c4664
15a4335c
235708c3
36644206
5f3c780c
a0370380
001c8ccc
011cce0c
15c30001
68062dc3
075c4664
30c36ff3
0002341c
780c6ed2
0007af5c
2006a077
8cac20b7
1cc301c3
3dc325c3
01334664
a037780c
0cc38ccc
2dc315c3
46643ac3
c828301c
0001311c
335c6c0c
08c315c4
420621d7
00073664
002ba4dc
ce50301c
0001311c
42724c0c
02734c0f
740c78af
71a4275c
435c4037
06c30e64
2cc32806
46643ac3
7084475c
05e454c3
002a04dc
6ff3675c
341c36c3
60070008
002a32dc
10f8301c
0000311c
8c0c6c0c
20060217
31c321c3
d0c34664
c828301c
0001311c
335c6c0c
1cc315a4
42171a84
49c33664
a406702b
05546027
6047a606
a8060254
10f8301c
0000311c
8c0c6c0c
200605c3
31c321c3
80c34664
6ff3175c
341c31c3
401c0004
411cc828
29c30001
67d2c82b
435c700c
09c31984
00f32806
435c700c
09c31984
04001a3c
36c328c3
301c4664
311cc828
6c0c0001
1944435c
15c308c3
3bc32dc3
60c34664
501c6164
511c10f8
740c0000
08c38c4c
21c32006
466431c3
8c4c740c
20060dc3
31c321c3
c0074664
002392dc
41074593
001174dc
345c8197
c3c325c4
7024575c
9c3cc584
7c4c0080
611cc006
36830005
32dc6007
09c30009
31c3200b
0004341c
42dc6007
406b0021
648532c3
808962b7
401c8177
411cc828
601c0001
bf0022b8
10c30157
0e942047
a21ca7c3
700c1ea0
335c540c
023c0904
4f5c01c0
14c300a1
a7c30173
1a88a21c
540c700c
0904335c
01c0023c
2ac32026
0ac33664
301ca0cb
311c10f8
6c0c0000
05c38c0c
21c32006
466431c3
301c0277
311cc828
6c0c0001
15a4335c
82972cc3
25c32a00
59c33664
801c742b
60270020
801c0754
60470030
801c0354
b01c0040
b11c10f8
1bc30000
8c0c640c
200608c3
31c321c3
40c34664
c828601c
0001611c
335c780c
60f71984
22970cc3
59c324c3
a0d7742b
780c5664
1944535c
18c304c3
3ac34257
60c35664
0bc36164
ac4c600c
200604c3
31c321c3
1bc35664
8c4c640c
20060257
31c321c3
c0074664
0018b4dc
9000601c
0001611c
c828501c
0001511c
335c740c
06c315a4
438619c3
580b3664
341c32c3
60070002
001722dc
401c540c
7e0022b8
425c6c0c
033c0904
206601c0
46642dc3
0380af3c
335c740c
0ac315a4
22bc201c
42063d00
26c33664
0e3f423c
341c34c3
193c0001
6bd201c0
b86b740c
0006a037
00b70077
3dc38cec
00f34664
335c740c
02c315a4
3664586b
c828801c
0001811c
440c18c3
01c0963c
03803f3c
6037b86b
09c388cc
2dc313c3
466435c3
680c28c3
15c4335c
163c0ac3
420600c0
00073664
001244dc
700c48c3
0944335c
219707c3
fe40293c
201c3664
00071111
001232dc
323c22f3
3364ff70
f5dc6027
c1970010
25c4365c
075cc3c3
c0847024
00809c3c
20067c4c
0005111c
60073183
000902dc
880b29c3
341c34c3
60070004
000fc2dc
65c3a86b
c2f7c485
01370889
c828401c
0001411c
22b8101c
0047bc80
a7c30e94
1ea0a21c
540c700c
0904335c
01c0023c
00814f5c
017314c3
a21ca7c3
700c1a88
335c540c
023c0904
202601c0
36642ac3
a0cb0ac3
10f8301c
0000311c
8c0c6c0c
200605c3
31c321c3
03374664
c828301c
0001311c
335c6c0c
2cc315a4
2a0082d7
366425c3
742b59c3
0020801c
07546027
0030801c
03546047
0040801c
10f8b01c
0000b11c
640c1bc3
08c38c0c
21c32006
466431c3
601c40c3
611cc828
780c0001
1984335c
0cc360f7
24c322d7
742b59c3
5664a0d7
535c780c
04c31944
431718c3
56643ac3
616460c3
600c0bc3
04c3ac4c
21c32006
566431c3
640c1bc3
03178c4c
21c32006
466431c3
7594c007
9000601c
0001611c
c828501c
0001511c
335c740c
06c315a4
438619c3
580b3664
341c32c3
60070002
540c5a54
22b8401c
6c0c7e00
0904425c
01c0033c
2dc32066
af3c4664
740c0380
15a4335c
201c0ac3
3d0022bc
36644206
423c26c3
34c30e3f
0001341c
01c0193c
740c6bd2
a037b86b
00770006
8cec00b7
46643dc3
740c00f3
15a4335c
586b02c3
801c3664
811cc828
18c30001
963c440c
3f3c01c0
b86b0380
88cc6037
13c309c3
35c32dc3
28c34664
335c680c
0ac315c4
00c0163c
36644206
48c30ef2
335c700c
07c320e4
293c2197
3664fe40
7777201c
00f30fd2
4444201c
201c0173
01133333
8888201c
0000211c
201c0073
02c32222
fc761296
08040f56
3f36f016
60c3e696
101c91c3
20800e40
205c2537
323c6fe3
7fe50106
f88c533c
323ca277
3364fff0
06356027
4407a5f2
0027e4dc
44070073
893c0b94
001c5080
011cbbbb
59c30000
2827055c
225702b3
893c2bd2
301c4d80
311caaaa
29c30000
26a7325c
365c0133
333c7004
321c02c7
89c301c8
365c8384
c3c37024
055c59c3
c08425c4
7044365c
0400133c
1c8424b7
d65c2377
301c7064
311cc828
6c0c0001
15a4335c
05800f3c
22bc401c
42063a00
165c3664
313c6fe3
7fe50206
f88c233c
03542047
10544007
433c784c
84370c8b
033c796c
03f70b0b
0b4b533c
001ca3b7
98001ea0
784c0193
0c0b533c
433ca437
83f70b8b
1a88501c
43b79a80
03542207
10544007
642c19c3
0004341c
301c6bd2
311cc828
6c0c0001
06c36eac
29c32609
265c3664
32c36ff3
0008341c
69d26337
833790cb
6e206497
a35764b7
a377b620
9000a01c
0001a11c
1258001c
02b71800
1ac0293c
649742f7
b01c6477
b11c8000
701c0001
80061000
501c8577
ba8022b8
1d13a237
04f70457
231c20c3
04350fff
1000401c
e4d784f7
acf2a557
0040d21c
0040c21c
70c304d7
b21cf805
a21c0040
101c0040
111cc828
640c0001
15a4335c
1cc30bc3
366427c3
c828201c
0001211c
335c680c
0ac315a4
27c31bc3
465c3664
34c36ff3
0002341c
32546007
ce50501c
0001511c
341c740c
6ed20004
c828001c
0001011c
2217600c
335c440c
023c0904
206601c0
201c01b3
211cc828
680c0001
500c8217
0904335c
01c0023c
45172146
501c3664
511cc828
740c0001
0006e037
00b70077
1bc38cec
65172ac3
23d74664
33542007
c828201c
0001211c
8217680c
335c500c
023c0904
208601c0
36644297
c828501c
0001511c
0f3c740c
00370580
0ac38ccc
05801f3c
37c34297
365c4664
60476fe3
796c1294
2000341c
740c6ed2
4026e037
40b74077
0dc38cec
2bc31ac3
46646297
00535bc3
65575ac3
12946007
ffc0d21c
ffc0c21c
401cb805
411cc828
700c0001
15a4335c
1cc305c3
36644806
001ce805
011cc828
600c0001
7064265c
00079f5c
06c38d0c
64971dc3
e0074664
101c1f54
111cc828
640c0001
21e4335c
245c49c3
df5c25a4
a0770007
501ce0b7
5f5c0100
00060066
20260137
01b72177
8e2c01f7
13c302c3
604642d7
44574664
49a064d7
d7844477
8557c784
a02554c3
0357a577
c1e410c3
fff160dc
40074417
301c3e54
6fa01000
54c38317
103435e4
221c2dc3
301c1000
311cc828
6c0c0001
00079f5c
06c38d0c
631712c3
401c4664
411cc828
700c0001
15a4335c
1cc30ac3
36644317
335c700c
19c321e4
25a4215c
0007df5c
0027af5c
80b78317
0100501c
00665f5c
01370006
21772026
01f701b7
02c38e2c
42d713c3
46646046
6ff3265c
341c32c3
265c0008
64f27044
4c2f38c3
831700b3
58c36a20
165c742f
08c37144
265c212f
400f7064
60ef6006
7124465c
365c810f
60476fe3
64070354
38c30c94
31c32cec
48c36572
a39770ef
313ca4d2
70ef0215
c828301c
0001311c
0fd203d7
335c6c0c
083c15a4
1f3c00c0
42060580
18c33664
617264ec
02d364ef
49c36c0c
25c4445c
58c34a00
065c342c
003771a4
0e64435c
0400023c
32c343d7
144f4664
627274ec
241774ef
10542007
4cec38c3
637232c3
70ef48c3
6ff3565c
341c35c3
64d20004
0185323c
365c70ef
62076fe3
64070354
29c30f94
341c682c
6ad20004
c828301c
0001311c
6eac6c0c
2a2906c3
365c3664
62076fe3
64070354
301c0b94
311cc828
6c0c0001
06c36e4c
366419c3
401c0693
411cc828
700c0001
1024335c
19c306c3
700c3664
06c3ae2c
29c32006
566431c3
09c3500c
25c4305c
f400401c
606c2e00
425c7112
001c15a4
011c8000
25800001
0c00201c
01f34664
0d944087
c828301c
0001311c
8e2c6c0c
29c32026
01215f5c
466435c3
fc761a96
08040f56
ff963016
12c351c3
c828301c
0001311c
335c6c0c
225c21e4
000625a4
8f8c0037
1ac0013c
23c312c3
466435c3
0c560196
00000804
315c3016
43c31629
1a546007
1609315c
61e78026
301c15b4
311cc828
2c0c0001
2449425c
02c7343c
01c8321c
1264415c
46642980
0b0d303c
433c33c4
04c3f88c
08040c56
3f36f016
70c3ec96
a264a1c3
826482c3
03c00f3c
42062006
0891bebc
02c00f3c
42062006
0891bebc
311c6c06
401c2200
411caaaa
8c0f0000
c828401c
0001411c
335c700c
012608c4
36642026
335c700c
01a608a4
36642026
6fa4975c
642c19c3
0004341c
a31c6dd2
0a540042
0034a31c
700c0754
07c36eac
29c32609
375c3664
63d26ee4
6d9460a7
0042a31c
301c0d94
311cc828
6c0c0001
15e4335c
c908001c
0010011c
a31c09d3
0d940034
c828301c
0001311c
335c6c0c
001c15e4
011cc930
07f30010
002ba31c
301c0d94
311cc828
6c0c0001
15e4335c
c958001c
0010011c
a31c0613
0d940025
c828301c
0001311c
335c6c0c
001c15e4
011cc978
04330010
0051a31c
301c0d94
311cc828
6c0c0001
15e4335c
c998001c
0010011c
a31c0253
04540026
002aa31c
301c0d94
311cc828
6c0c0001
15e4335c
c9a8001c
0010011c
301c3664
311cc828
6c0c0001
0624335c
8000001c
0001011c
28c31ac3
02f33664
311c6786
401c4105
411cab32
8c0f0000
c828301c
0001311c
8fec6c0c
101c07c3
111c8000
2ac30001
466438c3
ce54301c
0001311c
2c0f2006
6f84375c
900d201c
0000211c
34e442c3
19c3f894
341c642c
6bd20004
c828301c
0001311c
6eac6c0c
262907c3
366429c3
7184375c
a4dc6007
5c4c002d
1000241c
40074177
401c6d54
475c5aa5
875c6fc7
301c7007
311cc828
6c0c0001
07c36e6c
366419c3
30c340c3
2222361c
0b0d333c
633c7fe5
031cf88c
09541111
031cc8f2
05547777
031ca046
3f945555
ce54301c
0001311c
2c0f2006
ce58301c
0001311c
4c0d4006
c828301c
0001311c
6e0c6c0c
19c307c3
c5f23664
431ca026
25945555
6ee4375c
025460a7
301c6ef2
311cc828
6c0c0001
15e4335c
c9b8001c
0010011c
01333664
311c6786
201c4105
211cabf7
4c0f0000
c828301c
0001311c
6e8c6c0c
19c307c3
a0263664
c828301c
0001311c
6dec6c0c
19c307c3
366424c3
301c4d13
7d800e40
4f5c6277
34c300a1
0051a31c
60260294
c264c3c3
68f23cc3
002aa31c
a31c0554
d4dc0026
40060013
6f67275c
c828301c
0001311c
501c6c0c
511c9000
435c0001
05c315a4
cc24301c
0010311c
43862c0c
153c4664
053c00c0
3cc301c0
85c36ad2
a0c322b7
0033b55c
d01cb40b
01130000
22b7d5c3
b55ca0c3
b40b0033
353c8cc3
60070024
601c5f54
611cc828
580c0001
22b8401c
6c0c7e00
0904425c
01c0033c
42572146
780c4664
15a4335c
03c00f3c
22bc201c
42063d00
353c3664
101c0014
111ccc28
6fd20010
440c780c
0007bf5c
80778006
8cec80b7
12c30006
62572ac3
01134664
335c780c
0ac315a4
2bc3240c
501c3664
511cc828
540c0001
03c03f3c
88cc6037
13c30ac3
3bc34257
740c4664
15c4335c
03c00f3c
42062297
00073664
1cc32d94
740c28d2
0944335c
19c307c3
031328c3
335c740c
07c320e4
2dc319c3
301c0353
311cc828
201c0001
211ccc24
4cc30010
6c0c8ad2
0944335c
19c307c3
3664480c
01d340c3
335c6c0c
07c320e4
480c19c3
40c33664
1cc30753
5e542007
38c39fe6
323c4c89
7fe50036
66f27f32
04544027
2b944047
68d20133
ce50301c
0001311c
42724c0c
18c34c0f
60276489
301c0894
311cce50
4c0c0001
4c0f4072
648918c3
08946047
ce50301c
0001311c
41724c0c
301c4c0f
311cc828
6c0c0001
04a4335c
101c07c3
36642222
26948007
6ee4075c
00a703d2
301c1894
311cc828
4cc30001
6c0c89d2
15e4335c
c9dc001c
0010011c
6c0c0113
15e4335c
c9f4001c
0010011c
3fb33664
311c6786
101c4105
111cab53
2c0f0000
375c3e93
63d26ee4
249460a7
64f76006
22e0401c
0c0c7e00
64d70093
64f76025
30e464d7
301cfb14
311cc828
2cc30001
6c0c49d2
15e4335c
ca0c001c
0010011c
6c0cfad3
15e4335c
ca20001c
0010011c
6786f9d3
4105311c
abcc401c
0000411c
38738c0f
02b63a3c
233c7fe5
3a3cf88c
7fe50256
4bf27f32
a31c6af2
0a540042
a31c53c3
54dc0034
00930010
4d80693c
693c4af2
67f25080
02c7383c
01c8321c
d18049c3
38ef2006
ce0c301c
0001311c
980f8c8c
41f74c4c
2cac582f
4c6c384f
2d4c590f
4c0b392f
341c32c3
64f20001
0034a31c
24060794
7d6c38ef
0b0b233c
7c4c0093
0b8b233c
301c4237
311cce0c
4c0b0001
341c32c3
66d20004
64d26217
617278ec
78ec0073
78ef6272
115c19c3
908025c4
ce0cc01c
0001c11c
c828801c
0001811c
680c28c3
15a4335c
14c30cc3
36644806
0400d43c
8c0b3cc3
541c54c3
a0070004
000892dc
440c18c3
22b8301c
61377d80
425c6c0c
033c0904
206601c0
46644257
03c0bf3c
22bc401c
81b79e00
640c18c3
15a4335c
14c30bc3
36644206
02c05f3c
680c28c3
01804c3c
15a4335c
14c305c3
36644206
640c18c3
1584335c
220604c3
28c33664
bf5c680c
8ccc0007
1bc30cc3
68064257
48c34664
bf5c700c
8ccc0007
1bc30dc3
61d74257
18c34664
335c640c
0bc315c4
420615c3
00073664
42175794
29544007
1258301c
48c3bd80
2117700c
335c440c
023c0904
208601c0
366425c3
335c700c
0bc315a4
42062197
700c3664
0007bf5c
0dc38ccc
25c31bc3
466461d7
680c28c3
15a4335c
00c0063c
42061bc3
01d33664
700c48c3
71a4175c
435c2037
0dc30e64
421721d7
466432c3
a026184f
2cc303d3
48c3a8af
175c700c
203771a4
0e64435c
28060cc3
61d72dc3
784c4664
0c9430e4
640c18c3
71a4275c
435c4037
0dc30e64
25c321d7
a046fc13
c828301c
0001311c
335c6c0c
07c32124
1c80193c
366429c3
a02760c3
301c1f94
311c8000
ac0f0001
02b63a3c
7f327fe5
a31c64f2
27940025
201c69d2
211caaaa
19c30000
26a7215c
401c03d3
411cbbbb
39c30000
2827435c
a04702d3
3a3c1494
7fe502b6
64f27f32
0025a31c
275c0c94
49f27184
39c365d2
26a7235c
49c30093
2827345c
4006c5d2
215c19c3
375c246d
60077184
7c4c2494
1000341c
600760f7
a31c1e94
04540025
002ba31c
301c0b94
311cc828
6c0c0001
07c36e4c
366419c3
301c01d3
311cc828
6c0c0001
07c30e30
00613f5c
29c313c3
866431c3
175c2006
a0277187
301c1394
311cc828
c7f20001
6f2c6c0c
19c307c3
05d34a66
6f2c6c0c
19c307c3
00f4201c
a04704f3
375c2694
63d26ee4
0e9460a7
24f72006
22e0201c
4c0c7d00
64d70093
64f76025
32e464d7
301cfb14
311cc828
c8f20001
6f2c6c0c
19c307c3
00cc201c
6c0c00f3
07c36f2c
201c19c3
366400f6
fc761496
08040f56
0736f016
a0c3f896
315c71c3
20060564
1000111c
401c3183
411cf000
63d20000
0c24475c
341c7c2c
6bd20004
c828301c
0001311c
6eac6c0c
3e090ac3
366427c3
cc2c301c
0010311c
201c6c0c
211cccaa
4c0f0000
921c93c3
84c3c010
f000201c
601c8283
611cc828
780c0001
15a4335c
18c309c3
0ff8201c
780c3664
fff4243c
15a4335c
050019c3
4d40173c
36644c06
235c780c
573c21e4
175c1ac0
7c6c25a4
321c7112
6037d000
60776026
60b76006
01c38a0c
25c312c3
46646406
235c780c
175c21e4
7c6c25a4
321c7112
6037d000
00279f5c
1000301c
301c60b7
3f5c0100
60060066
60266137
60066177
61f761b7
01c38a2c
25c312c3
46646046
335c780c
275c21e4
8f5c25a4
20260007
20062077
8e0c20b7
13c302c3
640625c3
780c4664
21e4335c
25a4275c
00078f5c
00279f5c
1000101c
101c20b7
1f5c0100
20060066
20262137
20062177
21f721b7
02c38e2c
25c313c3
46646046
235c780c
175c21e4
7c6c25a4
321c7112
6037d000
60776026
60b76006
01c38a0c
25c312c3
46646406
341c7c2c
67d20004
6eac780c
3e290ac3
366427c3
08960006
0f56e076
00000804
43c33016
2476135c
2486235c
c828301c
0001311c
ae2c6c0c
24c32006
566431c3
08040c56
0136f016
50c3fe96
72c341c3
c21783c3
01212f5c
301c4077
311cc800
6c0c0001
23946007
311c6286
6c0c4105
0100341c
1b946007
6ee4305c
60a763d2
301c0e94
311cc828
6c0c0001
15e4335c
ca34001c
0010011c
01333664
311c6786
201c4105
211cab31
4c0f0000
02c7343c
335c7980
341c0f24
201c0001
211cc828
68d20001
2f5c680c
2f5c0021
8dcc0005
680c00f3
00212f5c
00052f5c
05c38dac
28c317c3
466436c3
80760296
08040f56
42c31016
6ee4305c
60a764d2
000a64dc
c800301c
0001311c
6ad26c0c
c828301c
0001311c
335c6c0c
000607e4
431c3664
62dc00f6
431c0008
11b400f6
5c548a67
05b48a67
f4dc8467
03530008
00cc431c
431c6b54
74dc00f4
0b530008
00fa431c
431c2754
05b400fa
00f9431c
02937c94
00fb431c
431c2954
759400fc
301c0633
311cc828
6c0c0001
15e4335c
ca44001c
0010011c
301c0c13
311cc828
6c0c0001
15e4335c
ca64001c
0010011c
301c0a93
311cc828
6c0c0001
15e4335c
ca80001c
0010011c
301c0913
311cc828
6c0c0001
15e4335c
ca98001c
0010011c
301c0793
311cc828
6c0c0001
15e4335c
cab4001c
0010011c
301c0613
311cc828
6c0c0001
15e4335c
cac4001c
0010011c
301c0493
311cc828
6c0c0001
15e4335c
cae0001c
0010011c
301c0313
311cc828
6c0c0001
15e4335c
cb24001c
0010011c
301c0193
311cc828
6c0c0001
15e4335c
cb50001c
0010011c
00f33664
ab00451c
311c6786
8c0f4105
08040856
0336f016
70c3fe96
41c303c3
82c34264
101c8264
111c8000
640c0001
0001341c
375c69f2
66d26ee4
045460a7
0001831c
343c3894
618002c7
0e84635c
0e44235c
0e64535c
fff0323c
ffff101c
03ff111c
39e491c3
202505b4
53e431c3
48c32635
4e948007
6ee4075c
00a703d2
301c0f94
311cc828
6c0c0001
15e4335c
cb94001c
0010011c
20463664
67860793
4105311c
ab4c201c
0000211c
60464c0f
06536077
c44c8489
a48c446c
02c7343c
315c2180
36e40e84
315c2594
32e40e44
315c2194
35e40e64
301c1d94
311cc828
6c0c0001
25c4405c
175c4a00
203771a4
0e64435c
0400023c
400615c3
466432c3
360330c3
0b0d333c
433c33c4
8077f88c
20260073
2f5c2077
02c30021
c0760296
08040f56
40c31016
0e240116
0014051c
80560f24
211c4246
680b4105
60723364
71cc680e
0004341c
19546007
c828301c
0001311c
6eac6c0c
145c04c3
243c0231
36640340
0704345c
0004341c
301c68d2
311c0600
4c0c4130
4c0f4072
311c6c06
40062200
00044c0f
321c0004
4c0c0420
48064c0c
00044c0f
00040004
f7de7a9c
08560013
00000804
02641016
436441c3
10540047
06b40047
00270dd2
000c34dc
00870133
00872d54
00a70d14
000bb4dc
201c0a13
211c0610
680c4130
159b303c
301c1613
311c0610
4c0c4130
213c2046
4c0f159b
111c2b86
201c4020
211c00b8
00664138
016f013c
6472680c
027f323c
311c6c86
03c34020
f49410e4
101c1273
111c0610
640c4130
323c4046
640f159b
311c6186
0c0e4020
211c4306
680c4138
680f6472
311c61c6
0c0e4020
680c4085
680f6472
311c6286
0c0e4020
680c4185
680f6472
311c62c6
0c0e4020
0cf34085
0610101c
4130111c
4046640c
159b323c
343c640f
6bd20014
311c6b86
40664020
201c4c0e
211c00b8
01334138
311c6186
00864020
43060c0e
4138211c
6472680c
343c680f
6bd20024
311c6bc6
40664020
201c4c0e
211c00bc
01334138
311c61c6
00864020
43860c0e
4138211c
6472680c
343c680f
6bd20044
311c6c46
40664020
201c4c0e
211c00c4
01334138
311c6286
00864020
45060c0e
4138211c
6472680c
343c680f
6bd20084
311c6c06
40664020
201c4c0e
211c00c0
01334138
311c62c6
00864020
45860c0e
4138211c
6472680c
0856680f
00000804
3f36f016
62c350c3
801cb3c3
78c30000
c828a01c
0001a11c
0034d01c
4105d11c
c01c9dc3
c11c003c
74cc4105
111c2006
31830010
1c546007
6ee4355c
60277fe5
1ac317b4
335c640c
07c30824
366415c3
44f228c3
0001801c
355c0293
101c6f84
111c900d
21c30000
f89432e4
355c0153
101c6f84
111c900d
21c30000
f89432e4
640c1dc3
a000341c
39c37cd2
6c0c4c0c
5fff101c
ffff111c
19c33183
241c640f
492700ff
49e70654
48a71254
03b32894
8000101c
0001111c
6f47155c
ab4f301c
0000311c
680f2cc3
0333e026
9000101c
0001111c
6f47155c
ab49301c
0000311c
680f2cc3
0173e006
6f84355c
900d101c
0000111c
32e421c3
05d3f894
0554ca27
0354c4c7
1e94c547
341c744c
60071000
1ac31994
335c640c
001c15a4
011cc830
155c0001
201c6f44
366405dc
05dc201c
6f67255c
900d301c
0000311c
6f87355c
1ac3eeb3
8d2c640c
16c305c3
1000201c
46643bc3
6006ed73
7187355c
0f56fc76
00000804
0336f016
90c3fe96
1264c257
23642077
73c34037
21c37364
6b5448c7
28c731c3
23c31cb4
02dc66e7
12c3000a
08b446e7
26a731c3
66c73e54
000da4dc
20570993
486721c3
000a12dc
288731c3
000a12dc
d4dc6707
11f3000c
21c32057
02dc4aa7
31c3000a
0db42aa7
6a6723c3
000b12dc
4a6712c3
000845dc
94dc2907
1193000b
32c34057
02dc6b47
12c30009
05544ea7
d4dc2ae7
1393000a
323c4017
798002c7
0f24335c
0020341c
2c946007
01936e26
323c4017
798002c7
0f24335c
0020341c
20946007
365c6626
1f5c2445
165c0001
11b3244d
323c4017
798002c7
0f24335c
0020341c
3f5c6fd2
365c0001
0ff32455
313c2017
798002c7
0f24335c
0020341c
301c6bd2
311cc828
6c0c0001
16c36f2c
00f9201c
305c0413
503c6e29
60675680
56c30254
c828801c
0001811c
4c0c38c3
02c7373c
01c8321c
1264425c
358009c3
466425c3
18c30ad2
6f2c640c
16c309c3
00fb201c
0e533664
323c4017
798002c7
0f87735c
60170893
24d6365c
165c2026
07b3246d
265c4006
0733246d
1221301c
2496365c
20260693
245d165c
40060613
245d265c
60260593
2465365c
20460513
2465165c
2f5c0493
265c0021
3f5c24b5
365c0001
765c24bd
301c24c6
311cc828
6c0c0001
13c4335c
366416c3
301c0213
311cc828
4c0c0001
313c2017
321c02c7
225c01c8
19801584
26642586
c828301c
0001311c
8e2c6c0c
200609c3
31c326c3
29c34664
6ee4025c
025400a7
301c0ef2
311cc828
6c0c0001
15e4335c
cba8001c
0010011c
01533664
21c32057
ab00251c
67864077
4105311c
02964c0f
0f56c076
00000804
1f36f016
70c3ff96
c82cc01c
0001c11c
611cc686
b01c4105
b11cc828
a01c0001
a11c003c
901c4105
911c0060
801c2200
811c0480
2cc32200
4dd24809
0e240116
0000041c
80560f24
6ee4375c
03946087
08d43cbc
341c780c
6007a000
780ced54
00ff341c
12946947
abaa201c
0000211c
4c0f3ac3
39c34006
28c34c0f
680c680c
00040004
8d9c0004
780cf7db
53c36037
5fff201c
ffff211c
780c5283
780f3283
680c2bc3
220b253c
07c38fac
00013f5c
353c13c3
4664808c
0196f7f3
0f56f876
00000804
0336f016
50c3fc96
20b71264
40772364
936493c3
6e29205c
0014323c
5680703c
703c63d2
60970340
88e743c3
002962dc
68e713c3
41c34fb4
a2dc26e7
34c30011
2ab486e7
666713c3
000c32dc
266741c3
34c31ab4
82dc8547
13c30008
0ab46547
24a741c3
000812dc
64c734c3
002aa4dc
80970ff3
256714c3
34c37b54
14dc6627
1233002a
14c38097
12dc26a7
86a7000e
000cc5dc
20970d33
684731c3
41c36954
0eb42847
872734c3
001812dc
472723c3
000ce0dc
882743c3
002844dc
20970fd3
488721c3
000b79dc
88c741c3
0027a4dc
209717d3
6aa731c3
000ad2dc
2aa741c3
34c323b4
d2dc8a07
13c30014
0eb46a07
294741c3
001362dc
696734c3
0015b2dc
290714c3
0025e4dc
609712b3
8a6743c3
0008c2dc
4a6723c3
0009a5dc
8a2743c3
002504dc
20973573
6b4731c3
000902dc
2b4741c3
34c30db4
92dc8ae7
13c30008
70dc6ae7
2b07001b
0023c4dc
40970bd3
6e4732c3
12c32b54
79542ea7
6e2732c3
002304dc
153c0333
40675680
17c30254
2493375c
1221331c
001bd2dc
6fa7155c
255c4097
401c6f07
411cc828
700c0001
05c36d6c
61063053
2200311c
23644c0b
4c0e4972
2449175c
61062077
2200311c
23644c0b
4c0e4972
c828301c
0001311c
8f8c6c0c
205705c3
602627c3
05c30593
40572006
084304bc
b2dc0007
301c001f
311cc828
00470001
6c0c0894
05c36f2c
201c17c3
00f300fb
6f2c6c0c
17c305c3
00fc201c
3cb33664
03944067
5680753c
c828301c
0001311c
8f8c6c0c
205705c3
604627c3
3ab34664
11944067
5680753c
355c01d3
6bd26ee4
095460a7
311c6786
101c4105
111cabf3
22d30000
c828301c
0001311c
e0376c0c
0404435c
2f5c05c3
12c30041
23c36057
466439c3
601c3653
611cc828
580c0001
2449475c
02c7343c
01c8321c
1264425c
3d8005c3
466427c3
25940007
2449175c
02c7313c
235c7d80
40070f84
355c3654
223c6e29
606702c7
780c0b94
0730221c
1264335c
350005c3
5680253c
780c0133
01c8221c
1264335c
3d0005c3
366427c3
1b540007
6ee4055c
0b5400a7
311c6786
201c4105
211cabf5
00070000
001644dc
c828301c
0001311c
335c6c0c
001c15e4
011ccbc4
27b30010
c828301c
0001311c
e0376c0c
0404435c
26e605c3
23c36057
466439c3
6ee4055c
0b5400a7
311c6786
101c4105
111cab37
00070000
000994dc
c828301c
0001311c
335c6c0c
001c15e4
011ccbdc
22b30010
311c6786
201c4105
211cabaa
4c0f0000
c828301c
0001311c
6f6c6c0c
366405c3
0e240116
0000041c
80560f24
311c6786
401c4105
411cabaa
8c0f0000
c82c301c
0001311c
2c0d2026
40672293
753c0394
801c5680
811cc828
48c30001
2057700c
02c7413c
1c80243c
1264335c
3d0005c3
366427c3
6f5c00f7
393c0061
60070014
c0071654
38c31494
7e004c0c
0e44135c
15c4425c
cc30301c
0010311c
275c0c0c
250025c4
46644806
c02602d2
8000301c
0001311c
8c0f8026
1394c007
6ee4055c
00a704d2
000c54dc
c828301c
0001311c
335c6c0c
001c15e4
011ccbf4
14b30010
74dcc027
055c000c
0ad26ee4
311c6786
101c4105
111cabcc
00a70000
301c0d94
311cc828
6c0c0001
15e4335c
cc04001c
0010011c
2c0f1153
201c1593
750022b8
60974c0c
6f07355c
c828401c
0001411c
6d6c700c
12c305c3
700c3664
05c36ecc
00414f5c
4f5c14c3
24c30021
12333664
c828601c
0001611c
101c580c
748022b8
425c6c0c
033c0904
308601c0
1258301c
46645580
1259401c
2c097600
241c21c3
40070004
74cc2754
211c4006
32830008
678669d2
4105311c
abcc401c
0000411c
301c0cf3
311cc828
6c0c0001
21e4335c
055c8eec
201c50e4
35001260
60264006
67864664
4105311c
abbb401c
0000411c
780c09f3
21e4335c
055c8eec
301c50e4
35801260
466432c3
311c6786
401c4105
411cabdd
07930000
6ee4055c
00a703d2
401c1694
411cc828
700c0001
15e4335c
cc14001c
0010011c
700c3664
15e4335c
cf30001c
0001011c
04733664
c828301c
0001311c
335c6c0c
001c15a4
011c8000
101c0001
111ccf30
46060001
67863664
4105311c
abaa201c
0000211c
01334c0f
311c6786
401c4105
411cabf3
8c0f0000
c0760496
08040f56
1f36f016
60c3ec96
72c3a1c3
60f73264
6ee4305c
08946047
211c4106
680b2200
feff341c
3a3c680e
9d8002c7
0e44045c
fff0303c
05dc7fa7
545c000c
453c0f24
40d70204
361c32c3
33c40002
f88cc33c
3cc383d2
800767f2
80d71094
202714c3
301c0c54
311cc828
6c0c0001
06c36f2c
201c17c3
153300f9
0400903c
0014353c
c828501c
0001511c
0100bf3c
21546007
821c86c3
540c1258
22b8401c
6c0c7a00
0904425c
01c0033c
28c32086
740c4664
175c09c3
408025c4
80378806
00770026
8cec00b7
12c309c3
38c32bc3
01734664
335c740c
0bc315a4
475c29c3
2a0025c4
36644806
00833f5c
5aa5331c
784c6594
2000341c
24946007
311c6286
6c0c4105
0100341c
1c946007
28f21cc3
4006796c
4000211c
60073283
501c1394
511cc828
540c0001
02c73a3c
01c8321c
1264425c
3d8006c3
466427c3
740c03d2
301c0853
311cc828
6c0c0001
4f5ce037
4f5c0061
8f0c0025
1ac306c3
01002f3c
466439c3
30c300d7
0002341c
67866ad2
4105311c
abaa101c
0000111c
05132c0f
d028301c
0001311c
47d24c09
6ee4365c
039460a7
086136bc
311c6786
001c4105
011cabaa
0c0f0000
c828301c
0001311c
6f6c6c0c
366406c3
301c0173
311cc828
6c0c0001
06c36f2c
446617c3
14963664
0f56f876
00000804
f896f016
311c6486
00464110
201c0c0e
211cd800
325c0001
101c6f84
111cbaad
01c30000
4a9430e4
6fa4625c
6f44725c
6f24025c
6f64325c
101c20c3
2183f000
21807fe5
f000301c
12e41383
10e40394
301c1494
311cc828
4c0c0001
ce0c301c
0001311c
6c4cac8c
890cc037
d800001c
0001011c
466425c3
d800301c
0001311c
6f64235c
25a4165c
6f24035c
e0770037
201c40b7
2f5c0100
60060066
00266137
61b70177
01c361f7
d69c101c
0010111c
1ac0263c
72bc6046
301c08a2
311cd800
101c0001
111c900d
135c0000
08966f87
08040f56
301c4006
311ccef4
4c0f0001
ce60301c
0001311c
201c4c0f
211ccf08
301c0001
311ccf00
280c0001
08042c0f
cf0c301c
0001311c
4c0f4006
ced4301c
0001311c
36646c0c
00000804
cef4201c
0001211c
cef8301c
0001311c
2c0f280c
ce60201c
0001211c
cefc301c
0001311c
2c0f280c
cf00201c
0001211c
cf04301c
0001311c
2c0f280c
00000804
cef8201c
0001211c
cef4301c
0001311c
2c0f280c
cefc201c
0001211c
ce60301c
0001311c
2c0f280c
cf04201c
0001211c
cf00301c
0001311c
2c0f280c
00000804
cf0c201c
0001211c
cf10301c
0001311c
2c0f280c
c828301c
0001311c
335c6c0c
36640504
00000804
cf10201c
0001211c
cf0c301c
0001311c
2c0f280c
c828301c
0001311c
335c6c0c
36640524
00000804
00734006
00254980
7df26008
118b323c
033c6d00
080403f4
30c3ff96
60373064
00012f5c
0604323c
04946807
46924017
323c00f3
67e707f4
40170494
40374672
00013f5c
019603c3
00000804
ff963016
306430c3
501c6037
511ccf0c
740c0001
15546007
ced8301c
0001311c
301c8c0c
311cc828
6c0c0001
05a4335c
00011f5c
366401c3
40064664
03b3540f
ced1301c
0001311c
20176c08
32e421c3
60260494
0233740f
ce84201c
0001211c
6025680c
301c680f
311cced8
6c0c0001
00011f5c
366401c3
0c560196
00000804
30c3ff96
60373064
cef4301c
0001311c
60076c0c
201c1294
211ccf00
680c0001
00011f5c
00df133c
201c680f
211cce60
680c0001
680f7fe5
08040196
cf08301c
0001311c
301c0c0f
311cced4
201c0001
211c51a4
4c0f0010
ced8301c
0001311c
5388201c
0010211c
08044c0f
51c37016
401c62c3
411cc828
700c0001
0604335c
700c3664
06e4335c
16c305c3
0e563664
00000804
301c7016
311ccecc
8c0c0001
c828601c
0001611c
ced0501c
0001511c
780c00f3
1504335c
36641409
80079fe5
0e56f9d4
00000804
ff963016
401c50c3
411cc828
700c0001
0644335c
01333664
700ca025
1504335c
00012f5c
366402c3
60377408
019676f2
08040c56
fe967016
cf14401c
0001411c
500d4026
702d6466
0200303c
2f5c6077
504d0021
706d6b26
d08dc006
c828501c
0001511c
335c740c
043c0584
36640010
0200303c
2f5c6037
508d0001
cec8301c
0001311c
50ad4c09
740cd0cd
0664335c
366404c3
0e560296
00000804
fe967016
cf14401c
0001411c
500d4026
702d6466
0200303c
2f5c6077
504d0021
706d69c6
d08dc006
c828501c
0001511c
335c740c
043c0584
36640010
0200303c
2f5c6037
508d0001
cec8301c
0001311c
50ad4c09
740cd0cd
0664335c
366404c3
0e560296
00000804
0136f016
80c3fb96
cec8301c
0001311c
0c0d01a6
cecc301c
0001311c
2c0f2006
ced0301c
0001311c
4c0d4006
ced1301c
0001311c
8c0d8466
cef0101c
0001111c
301c440c
311ccc34
0c0c0010
24e440c3
323c0494
640ffff0
cedc701c
0001711c
cef0301c
0001311c
6fa06c0c
6007a066
7fe574f4
cf14401c
0001411c
308d2fc6
6007a086
7fe56a54
50ad44a6
6007a0a6
233c6454
7c49fff0
1c0503c3
301c0137
311ccecc
1f5c0001
2c0f0081
70cd6406
4007a0c6
623c5254
301cfff0
311cc828
6c0c0001
05a4335c
36641c69
ced0301c
0001311c
08060c0d
a0e610ed
3d54c007
fff0263c
31c33c89
60f77c05
cec8301c
0001311c
00610f5c
25a60c0d
a106310d
2b544007
301c5fe5
311cced1
1ca90001
24660c0d
a126312d
1f544007
fff0323c
514d49c6
6007a146
7fe51854
116d0626
6007a166
29c61254
a186318d
0d546027
cf14301c
0001311c
8dad8446
0dcd0406
2ded2606
a2060e0d
cf14401c
0001411c
500d4026
0200053c
1f5c00b7
302d0041
0200383c
0f5c6077
104d0021
306d2b26
4006a025
601c52a1
611cc828
780c0001
0584335c
0010043c
103c3664
20370200
00012f5c
253c52a1
301c0010
311ccec8
0c090001
6a001121
2c2d2006
335c780c
04c30664
05963664
0f568076
00000804
3f36f016
a0c3fe96
501c2037
511cce84
00060001
301c140f
311ccec8
21a60001
301c2c0d
311ccecc
0c0f0001
ced0301c
0001311c
4c0d4006
ced1301c
0001311c
0c0d0466
c828401c
0001411c
335c700c
366404e4
335c700c
36640544
0000901c
d01cdfe6
d11ccef0
74c30001
c5c3b4c3
cedc201c
0001211c
440f1dc3
035c7c0c
06641524
326430c3
04546027
f7946067
2bc32b33
035c680c
06641524
506450c3
0e04353c
12dc6007
0bc3000c
035c600c
06641524
406440c3
0e04343c
52dc6007
343c000b
933cfe00
96e40ff4
2bc30694
335c680c
00b30564
600c0bc3
0544335c
7c0c3664
1524035c
80c30664
383c8064
60070e04
000992dc
0ff4243c
0ff4353c
383c4980
c9800ff4
fe00353c
00ff341c
ffe0433c
6b946007
035c7c0c
06641524
506450c3
0e04353c
7e546007
035c7c0c
06641524
406440c3
0e04343c
74546007
035c7c0c
06641524
303c0064
60070e04
353c6b54
4f000ff4
0ff4343c
313c2980
6c80118b
003f341c
03e46405
343c5d94
233cfe00
353c0ff4
341cfe00
333c00ff
898005f7
0ff4303c
0633cc80
035c7c0c
06641524
306430c3
341c6077
600700e0
831c4354
09940044
335c7c0c
2f5c05c4
02c30021
02b33664
0053831c
0dc31294
31c3200c
00212f5c
00df233c
001c600f
011ccc38
400c0010
031432e4
280f2dc3
30c30057
00ff341c
9fe5d980
cfd48027
680c2bc3
1524035c
20c30664
323c2064
60070e04
363c1154
6f00118b
003f341c
23e46405
7c0c0994
1524035c
30c30664
61a73264
69c30c54
335c7c0c
36640564
335c7c0c
09c306a4
e3733664
0053831c
7c0c0794
06c4335c
366409c3
831c0f33
6e940044
d800101c
0001111c
6f84315c
900d001c
0000011c
32e420c3
301cf494
311ccf08
4c0c0001
8000001c
0001011c
23e430c3
001c1394
011ccf00
600c0001
0cc36d20
001c600f
011c9000
301c0001
311ccf08
0c0f0001
201c0353
211ccf00
680c0001
9000001c
0001011c
2cc36c20
001c680f
011c8000
301c0001
311ccf08
0c0f0001
9000201c
0001211c
6f47215c
335c7c0c
366404e4
0051a31c
a31c0754
04540026
002aa31c
201c1094
211cd800
684c0001
1000341c
7c0c68f2
02c36d4c
280c2cc3
01933664
8d2c7c0c
d800001c
0001011c
3cc31ac3
60174c0c
7c0c4664
0684335c
366409c3
0042831c
69c30554
0006d313
301c0193
311ccf00
4c0c0001
cf08301c
0001311c
08a02c0c
fc760296
08040f56
fe961016
2f5c4006
40060036
111c2f86
640b4010
3f5c3364
3f5c0036
033c0033
0af20084
60064045
0200311c
24e443c3
0037f194
60060273
4010311c
23c36c0b
40372264
c828301c
0001311c
335c6c0c
4f5c1504
04c30001
2f5c3664
02c30001
08560296
00000804
0136f016
2006fc96
00561f5c
00661f5c
2f5c4626
301c007d
311cd800
335c0001
83c36e29
341c6ad2
801c0001
811cd834
63f20001
0534821c
ce5c301c
0001311c
20072c09
001414dc
325c28c3
331c2584
0d9400f1
c828301c
0001311c
335c6c0c
001c15e4
011ccc3c
01f30010
00f2331c
301c0d94
311cc828
6c0c0001
15e4335c
cc5c001c
0010011c
401c3664
411cc828
700c0001
15e4335c
cc78001c
0010011c
700c3664
15e4335c
cc98001c
0010011c
700c3664
15e4335c
ccb4001c
0010011c
301c3664
311cd800
335c0001
65f26ee4
335c700c
366414c4
c828401c
0001411c
335c700c
001c15e4
011cccb8
36640010
335c700c
001c15e4
011cccdc
36640010
335c700c
001c15e4
011ccd08
36640010
335c700c
001c15e4
011ccd34
36640010
335c700c
001c15e4
011ccd6c
36640010
d800301c
0001311c
341c6d6c
60070001
700c3154
15e4335c
cda4001c
0010011c
700c3664
15e4335c
cdc4001c
0010011c
700c3664
15e4335c
cdec001c
0010011c
700c3664
15e4335c
ce14001c
0010011c
700c3664
15e4335c
ce44001c
0010011c
700c3664
15e4335c
ce78001c
0010011c
401c3664
411cc828
700c0001
15e4335c
cea0001c
0010011c
700c3664
15e4335c
cec4001c
0010011c
700c3664
15e4335c
cee8001c
0010011c
700c3664
15e4335c
cef8001c
0010011c
18c33664
2459315c
5e946027
335c700c
001c15e4
011ccf0c
36640010
335c700c
001c15e4
011ccf28
36640010
335c700c
001c15e4
011ccf44
36640010
335c700c
001c15e4
011ccf5c
36640010
335c700c
001c15e4
011ccf74
36640010
335c700c
001c15e4
011ccfa4
36640010
d800301c
0001311c
6e29135c
341c31c3
69d20001
335c700c
001c15e4
011ccfcc
36640010
d800201c
0001211c
341c696c
60070001
125c1354
31c36e29
0002341c
301c6dd2
311cc828
6c0c0001
15e4335c
cfe4001c
0010011c
301c3664
311cc828
6c0c0001
15e4335c
ccb4001c
0010011c
301c3664
311cc828
6c0c0001
00078f5c
0764435c
d800001c
0001011c
00f01f3c
60064026
30c34664
60073264
000e94dc
00792f5c
fbf0123c
3f5c2077
60270021
46671335
46871154
48c70f54
46a70d54
46c70b54
49670954
47270754
4ae70554
4a670354
48c76894
48270b54
48470954
46a70754
49670554
4ae70354
301c0d94
311cc828
6c0c0001
15e4335c
cff8001c
0010011c
301c0193
311cc828
6c0c0001
15e4335c
d01c001c
0010011c
601c3664
611cc828
780c0001
00795f5c
00078f5c
0764435c
d800001c
0001011c
00a01f3c
35c34046
30c34664
60073264
000944dc
00793f5c
f4dc68c7
780c0008
15e4335c
d038001c
0010011c
780c3664
15e4335c
d060001c
0010011c
780c3664
00795f5c
00078f5c
0764435c
d800001c
0001011c
00c01f3c
35c34066
30c34664
60073264
14536a54
42944b47
c828701c
0001711c
335c7c0c
001c15e4
011cd078
36640010
5f5c7c0c
8f5c0079
435c0007
001c0764
011cd800
1f3c0001
408600a0
466435c3
326430c3
47946007
00536f5c
4394c0a7
335c7c0c
001c15e4
011cd090
36640010
5f5c7c0c
8f5c0079
435c0007
001c0764
011cd800
1f3c0001
26c300c0
466435c3
326430c3
27546007
46e70bf3
401c2494
411cc828
700c0001
15e4335c
d0ac001c
0010011c
700c3664
00795f5c
00078f5c
0764435c
d800001c
0001011c
00a01f3c
35c340c6
30c34664
65d23264
262607b3
007d1f5c
325c28c3
331c2493
14941221
00793f5c
03546847
0e946687
c828301c
0001311c
335c6c0c
001c15e4
011cd0e8
36640010
301c0433
311cd800
335c0001
69f26ee4
c828301c
0001311c
335c6c0c
366414c4
c828301c
0001311c
8fac6c0c
d800001c
0001011c
00791f5c
00532f5c
00633f5c
04964664
0f568076
00000804
401c3016
411cc828
501c0001
511cce5c
700c0001
0724335c
700c3664
15e4335c
d120001c
0010011c
60263664
fe53740d
08040c56
1f36f016
90c3f896
62c341c3
200683c3
00f61f5c
701ca006
711cc828
c01c0001
a01c0b00
a11c007c
b01c4010
b11c0000
a0254010
325c29c3
60076ee4
1ac31194
3364640b
00f63f5c
00f33f5c
0008341c
82dc6007
2bc3000e
700d680b
3cc301d3
305c0c0c
6ceb0b64
c2dc6007
101c000d
5ebc0200
100d08c6
335c7c0c
10091504
c0673664
000982dc
07b4c067
0f54c027
84dcc047
0e53000b
d2dcc0a7
c0a70008
000a30dc
e4dcc0c7
13d3000a
46275009
48273354
48473154
46872f54
46a72d54
46c72b54
46e72954
47072754
49672554
47272354
4a272154
44c71f54
45471d54
48671b54
48871954
49071754
4aa71554
45671354
44a71154
46670f54
4b470d54
48c70b54
4ae70954
48e70754
4a870554
4a670354
24977794
2459315c
0a546027
08544867
06544a87
04544ae7
64dc4a67
46270008
000832dc
02dc4827
48470008
46877d54
49677b54
47277954
7c0c7754
15e4335c
d138001c
0010011c
7c0c3664
0704335c
00073664
7c0c6994
15e4335c
d168001c
0010011c
70090293
1b946607
0034831c
831c0754
04540036
0039831c
7c0c1294
15e4335c
d1ac001c
0010011c
7c0c3664
15e4335c
d188001c
0010011c
07333664
123c5009
20f7fd00
00613f5c
61276177
2f5c04b4
033300a1
f9f0323c
3f5c60b7
60a70041
123c15b4
2077fa90
00212f5c
30090193
5a0521c3
3f5c4037
61b70001
06b460a7
00c12f5c
6006500d
7c0c0373
15e4335c
d1cc001c
0010011c
7c0c3664
15e4335c
d188001c
0010011c
a0253664
fffe101c
01ff111c
52e421c3
fff019dc
61376026
20060073
2f5c2137
02c30081
f8760896
08040f56
ff963016
d800301c
0001311c
6ee4335c
60076037
44bc2194
30c3082d
1f5c3264
21c30001
029469c7
42c34026
6b274264
80070354
44bc3b54
30c3082d
68a73264
80073594
44bc3394
30c3082d
04c33264
2d946a67
301c0533
0c0c0b00
0200101c
08c65ebc
326430c3
04e6233c
423c5fe5
6b27f88c
80070354
501c1954
140c0b00
0200101c
08c65ebc
326430c3
0e9468a7
140c8df2
0200101c
08c65ebc
326430c3
6a6704c3
00260494
00060053
0c560196
00000804
401c3016
411cc828
700c0001
20a4335c
700c3664
1d04335c
d800001c
0001011c
501c3664
700c0b00
1ce4335c
3664140c
335c700c
140c1d24
f3243664
08040c56
40c31016
8000301c
0001311c
2c0f2026
6ee4305c
11946087
0e240116
0014051c
80560f24
c828301c
0001311c
335c6c0c
04c30784
04f33664
1c946027
4006604c
8000211c
6ed23283
cf30301c
0001311c
135c2b26
301c0155
311c0254
43262020
62464c0e
4105311c
23644c0b
4c0e4072
60470153
301c0894
311c800c
4c0c4600
4c0f4f92
6e29345c
17546007
2724245c
245c46f2
49d250c4
07946047
ab00251c
311c6786
01134105
311c6786
201c4105
211cab10
4c0f0000
c828301c
0001311c
6fcc6c0c
366404c3
6ee4345c
08946087
0116f524
051c0e24
0f240000
08568056
00000804
301cfd96
311cc828
6c0c0001
0a64335c
20460fc3
301c3664
311c801c
201c4113
4c0e0100
08040396
50c33016
301c5264
311cd800
335c0001
60a76ee4
01162294
051c0e24
0f240014
301c8056
311cc828
6c0c0001
0784335c
401c3664
100c0b00
0200101c
08c65ebc
0abc0aa6
100c0861
0200101c
08c65ebc
326430c3
f0946aa7
301cadd2
311cc828
6c0c0001
15e4335c
d1e0001c
0010011c
301c3664
311cc828
6c0c0001
0744335c
301c3664
311cd800
335c0001
60a76ee4
f5240894
0e240116
0000051c
80560f24
08040c56
ff963016
501c40c3
511cc828
01330001
335c740c
2f5c1504
02c30001
80253664
60377009
019676f2
08040c56
0364ff96
311c6206
0c0e4001
311c6186
20264001
42862c0e
4001211c
3364680b
341c6037
7bd28000
00012f5c
019602c3
00000804
2037ff96
402744d2
00b30994
00013f5c
00d3600d
600e6017
60170073
0196600f
00000804
1f36f016
83c3a1c3
311c6386
101c4001
2c0e0141
4b544007
af7250c3
733c6026
c7c4800d
97a492c3
c828b01c
0001b11c
640c1bc3
0ac4335c
366405c3
626460c3
28c3a025
25544007
640c1bc3
0ac4335c
366405c3
400c303c
ff00341c
a02563a3
0001831c
1bc31635
335c640c
05c30ac4
40c33664
a0254264
680c2bc3
0ac4335c
366405c3
c00c303c
81ac343c
a02563a3
640c1bc3
0ae4335c
16c30ac3
366428c3
29c39c84
63d26b80
f873a784
0f56f876
00000804
311c6706
44064140
08044c0e
00000804
205c40c6
67866ee7
4105311c
ab10201c
0000211c
301c4c0f
311cc828
6c0c0001
36646fcc
00000804
211c4506
080f4105
8170201c
4600211c
0804080f
311c6006
101c4140
2c0f0300
311c6486
201c0080
211c0000
4c0f0800
101c6085
111c0000
2c0f0400
201c6105
211c0000
4c0f0800
101c6085
111c0000
2c0f0800
211c4286
60260080
301c680f
311c0084
20464105
680c2c0f
0001341c
42867dd2
0080211c
6007680c
0804fe15
226420c3
311c6286
6c0c4105
0100341c
14dc6007
6006000e
4140311c
111c2006
2c0f0040
3c544067
07b44067
0d544027
a4dc4047
0313000c
715440a7
4c1440a7
24dc40e7
1333000c
211c4006
21864130
6086280f
4130311c
2c0f2866
311c6006
680f00f0
40061633
4130211c
280f20c6
311c6086
29264130
20062c0f
00d0111c
4006280f
0020211c
4b064c0f
4600211c
2006680c
0400111c
7bd23183
400612b3
4130211c
680f6106
311c6086
28e64130
20062c0f
00b0111c
4006280f
0040211c
4b064c0f
4600211c
2006680c
2000111c
7bd23183
40860f33
4130211c
680f69e6
311c6006
20064130
0090111c
60062c0f
0060311c
4b06680f
4600211c
2006680c
0400111c
7bd23183
211c4b06
680c4600
111c2006
31832000
0ad37bd2
211c4006
68264130
6086680f
4130311c
2c0f21c6
111c2006
280f0010
211c4006
4c0f00e0
211c4686
680c4140
111c2006
31830004
4b067bd2
4600211c
2006680c
0400111c
7bd23183
211c4b06
680c4600
111c2006
31832000
05137bd2
311c6006
40264130
60854c0f
111c2006
2c0f00f0
4c0f49c6
211c4686
680c4140
111c2006
31830002
4b067bd2
4600211c
2006680c
0400111c
7bd23183
211c4b06
680c4600
111c2006
31832000
60867bd2
4140311c
211c4006
4c0f0040
00000804
ff963016
301c51c3
311cc828
6c0c0001
71a4205c
435c4037
013c0e64
101c1c80
400602e4
466432c3
2567055c
0c560196
00000804
0136f016
80c3ff96
000651c3
2587015c
1c80613c
c828701c
0001711c
215c7c0c
335c25e4
06c315a4
25c4415c
201c2a00
366402e8
08c37c0c
71a4005c
435c0037
06c30e64
02e4101c
32c34006
155c4664
21c32564
355402e4
355c5c0c
401c25c4
2e00e000
7112746c
15a4425c
258006c3
02e8201c
7c0c4664
005c08c3
003771a4
0e64435c
101c06c3
400602e4
466432c3
155c2006
255c246d
42c32564
0d5404e4
00f2001c
2587055c
335c7c0c
06c31584
02e8101c
00b33664
00f1101c
2587155c
80760196
08040f56
ff961016
31c3240c
411c8006
34830100
31c36cd2
211c4006
32830400
22546007
305c6026
03d36e25
411c8006
14830200
27d22037
305c6026
205c6e3d
00b36e47
00014f5c
6e3d405c
6e39205c
301c4bd2
311cc828
6c0c0001
09a4335c
6e44005c
01963664
08040856
24d2ff96
06942027
60090073
600b0093
600c0053
60176037
019603c3
00000804
00000804
0736f016
50c3ff96
72c301c3
8f5c43c3
c0260124
073538e4
04946047
38c3c086
c04662d2
4c54e007
400616c3
831c4037
13540001
65d238c3
0002831c
03331d94
180c923c
a3c36aa2
6017a923
9aa393c3
00079f5c
02134025
180c923c
a3c36ae2
6017a923
9aa393c3
00079f5c
00934045
4037540c
3fe54086
da942007
44f232c3
b580fda0
8027fa13
84d20e54
12548047
1f5c02d3
103c0001
201700df
20372832
fdd35fe5
103c2017
3032016f
5fc52037
4017fcf3
027f203c
fc534006
01960013
0f56e076
00000804
6232600b
7fe50004
fd947fe7
00000804
0336f016
30c3ff96
92c351c3
2c4c002c
243c8c0c
643c150b
34c3158b
833c3364
433c0010
34c3801b
711ce006
37830100
20946007
600674c3
8000311c
e6d27383
0f24355c
355c6872
301c0f27
311cc828
6c0c0001
00079f5c
0be4435c
36c328c3
e0074664
355c1254
68920f24
0f27355c
301c0193
311cc828
6c0c0001
435c4037
28c310c4
466436c3
c0760196
08040f56
40c33016
c828501c
0001511c
500c740c
1084335c
123c102c
3664150b
304c30c3
506c3183
31e412c3
0c56f294
00000804
20c31016
c828301c
0001311c
800c6c0c
0ae4335c
284c002c
158b243c
08563664
00000804
40c33016
c828501c
0001511c
400c740c
1084335c
123c004c
3664150b
702c10c3
740c1383
335c500c
106c0ae4
15a3b08c
158b223c
0c563664
00000804
313c200b
67d20014
8020301c
4113311c
4c0e4c06
0024313c
404b67d2
8028301c
4113311c
313c4c0e
66d20044
6186404c
4140311c
313c4c0f
66d20084
6206406c
4140311c
313c4c0f
66d20104
6286408c
4140311c
313c4c0f
69d20204
c828301c
0001311c
6c6c6c0c
366400ac
00000804
3f36f016
80c3f896
72c391c3
042b64d2
007301f7
21f724d7
c828501c
0001511c
00406f3c
0014d01c
4105d11c
0080cf3c
01c0bf3c
e037740c
0be4435c
16c301d7
60464086
40574664
240b323c
d200401c
0010411c
3a1da43c
600c0dc3
0100341c
18c36bd2
6e31115c
32c32ed2
411c8006
34832000
32c300d3
011c0006
30834000
43546007
e037740c
0be4435c
033c61d7
1cc30040
ffc02a3c
46646046
00331f5c
341c31c3
6047000f
60471a54
6bd205d4
27946027
60870193
60871a54
60a71474
03332094
335c740c
031310e4
335c740c
06c31104
27c318c3
02f33664
335c740c
01931124
335c740c
01131144
335c740c
00931164
335c740c
06c31184
00b33664
335c740c
366410a4
31c32057
011c0006
30830600
211c4006
42c30200
155434e4
61d72ac3
01f70980
800631c3
0800411c
60073483
740c8054
435ce037
1bc30be4
60464086
eef34664
c828301c
0001311c
335c6c0c
08c31064
0700193c
53ac49c3
08963664
0f56fc76
00000804
70c3f016
52c341c3
450c63c3
1004323c
10946007
341c750c
6cd20100
687232c3
f1ff101c
710f3183
241c550c
32a30e00
710c710f
0004341c
22946007
341c750c
60070004
301c1d54
311cc828
6c0c0001
15a4335c
0340043c
0340153c
36644186
32c3510c
710f6272
2006750c
0800111c
66d23183
311c6086
23a30800
750c510f
0008341c
352c6bd2
365c312f
63922684
2687365c
6372710c
750c710f
0010341c
554c6bd2
365c514f
64922684
2687365c
6472710c
750c710f
0020341c
756c6bd2
365c716f
65922684
2687365c
6572710c
750c710f
0040341c
358c6bd2
365c318f
66922684
2687365c
6672710c
750c710f
1000341c
560c6bd2
365c520f
6c922684
2687365c
6c72710c
750c710f
2000341c
762c6bd2
365c722f
6d922684
2687365c
6d72710c
750c710f
4000341c
364c6bd2
365c324f
6e922684
2687365c
6e72710c
355c710f
67320109
566c6bd2
365c526f
6f922684
2687365c
6f72710c
750c710f
111c2006
31830100
568c6bd2
365c528f
78922684
2687365c
7872710c
750c710f
111c2006
31831000
710c64d2
710f7c72
0101355c
60076732
542c1754
744c502f
346c704f
548c306f
74ac508f
34cc70af
54ec30cf
710c50ef
710f6772
2684365c
365c6792
245c2687
323c0484
6cf20014
0484355c
0001341c
32c367d2
345c6072
742b0487
245c702e
323c0484
60070024
355c1794
341c0484
60070002
155c1154
145c04c1
355c04c5
345c04c9
155c04cd
145c04d1
32c304d5
345c6172
245c0487
32c304a4
1000341c
355c6af2
341c04a4
65d21000
6c7232c3
04a7345c
04a4245c
341c32c3
6af22000
04a4355c
2000341c
32c365d2
345c6d72
245c04a7
323c0484
6af20044
0484355c
0004341c
32c365d2
345c6272
355c0487
341c0484
6ed20008
04e4255c
04e7245c
0504355c
0507345c
0484345c
345c6372
355c0487
20060484
4000111c
6ad23183
0524255c
0527245c
0484345c
345c7e72
245c0487
323c0484
6ef20104
0484355c
0010341c
355c69d2
345c0544
32c30547
345c6472
245c0487
323c0484
6ef20204
0484355c
0020341c
155c69d2
145c0564
32c30567
345c6572
245c0487
323c0484
6ef20404
0484355c
0040341c
355c69d2
345c0584
32c30587
345c6672
345c0487
67320481
18946007
0481355c
60076732
301c1354
311cc828
6c0c0001
15a4335c
0c00043c
0c00153c
36644206
0484345c
345c6772
245c0487
323c0484
60071004
355c1294
341c0484
6dd20100
0684155c
0687145c
06a4355c
06a7345c
687232c3
0487345c
0484245c
4004323c
355c6ef2
341c0484
69d20400
06c4155c
06c7145c
6a7232c3
0487345c
0484245c
8004323c
355c6ef2
341c0484
69d20800
06e4355c
06e7345c
6b7232c3
0487345c
0484345c
1000341c
19946007
0484355c
1000341c
13546007
c828301c
0001311c
335c6c0c
043c15a4
153c0e00
41860e00
345c3664
6c720484
0487345c
0484245c
341c32c3
60074000
355c1294
341c0484
6dd24000
0764155c
0767145c
0784355c
0787345c
6e7232c3
0487345c
0484245c
341c32c3
6df28000
0489355c
69d26732
07a4155c
07a7145c
6f7232c3
0487345c
0484245c
200632c3
0001111c
6df23183
0484355c
69d23183
07c4355c
07c7345c
707232c3
0487345c
0484245c
200632c3
0002111c
6df23183
0484355c
69d23183
07e4355c
07e7345c
717232c3
0487345c
0484245c
200632c3
0004111c
6df23183
0484355c
69d23183
0804355c
0807345c
727232c3
0487345c
0484245c
200632c3
0008111c
6df23183
0484355c
69d23183
0824355c
0827345c
737232c3
0487345c
0484245c
200632c3
0010111c
6df23183
0484355c
69d23183
0844355c
0847345c
747232c3
0487345c
0484245c
200632c3
0040111c
6df23183
0484355c
69d23183
0864355c
0867345c
767232c3
0487345c
0491345c
60076732
355c1894
67320491
13546007
c828301c
0001311c
335c6c0c
043c15a4
153c1100
43861100
345c3664
77720484
0487345c
0484245c
200632c3
0200111c
6df23183
0484355c
69d23183
0b24355c
0b27345c
797232c3
0487345c
0484245c
200632c3
1000111c
6df23183
0484355c
69d23183
0b44355c
0b47345c
7c7232c3
0487345c
0484245c
200632c3
2000111c
6df23183
0484355c
69d23183
0b64355c
0b67345c
7d7232c3
0487345c
04a4245c
0014323c
355c6ef2
341c04a4
69d20001
607232c3
04a7345c
05a4155c
05a7145c
04a4245c
0024323c
355c6ef2
341c04a4
69d20002
617232c3
04a7345c
05c4255c
05c7245c
04a4245c
0044323c
355c6ef2
341c04a4
69d20004
627232c3
04a7345c
05e4355c
05e7345c
04a4245c
2004323c
355c6cf2
341c04a4
67d20200
338f378c
697232c3
04a7345c
04a4245c
1004323c
355c6cf2
341c04a4
67d20100
73af77ac
687232c3
04a7345c
04a4245c
0084323c
355c6af2
341c04a4
65d20008
637232c3
04a7345c
04a4245c
0404323c
355c6ef2
341c04a4
69d20040
667232c3
04a7345c
0be4155c
0be7145c
04a4245c
0104323c
12946007
04a4355c
0010341c
32c36dd2
345c6472
255c04a7
245c0ba4
355c0ba7
345c0bc4
355c0bc7
20060484
0100111c
60073183
153c1754
7c2c1480
c828401c
0001411c
0080073c
700c69f2
15a4335c
36644386
5c2f4046
700c00b3
2104335c
0f563664
00000804
41c33016
313c200c
62070304
500c1d54
110b223c
323c31c3
600f111b
333c702c
402c0b0b
0b1b233c
702c402f
234b333c
133c12c3
202f235b
223c502c
31c3250b
251b323c
700c602f
0030341c
1e946207
313c304c
60070024
404c1954
0024323c
14946007
084b313c
085b233c
704c404f
208b333c
133c12c3
204f209b
223c504c
31c3250b
251b323c
200c604f
f004313c
500c68f2
220b223c
323c31c3
600f221b
306c606c
606f31a3
508c608c
608f32a3
32c3400c
35a3b00c
0b0b133c
313c32c3
600f0b1b
300c23c3
223c21a3
323c0b4b
600f0b5b
b00c23c3
223c25a3
323c0b8b
600f0b9b
300c23c3
223c21a3
323c0bcb
600f0bdb
25c3b02b
0001241c
0c0b133c
323c21a3
600f0c1b
300c23c3
223c21a3
323c0c4b
600f0c5b
b00c23c3
223c25a3
323c0c8b
600f0c9b
323c402c
60070014
702c3094
0001341c
2b546007
607232c3
23c3602f
21a3302c
084b223c
085b323c
23c3602f
25a3b02c
088b223c
089b323c
23c3602f
21a3302c
08cb123c
213c23c3
402f08db
333c702c
12c3190b
191b133c
502c202f
164b223c
323c31c3
602f165b
32c3402c
35a3b02c
0ecb133c
313c32c3
602f0edb
302c23c3
223c21a3
323c0f0b
602f0f1b
b02c23c3
223c25a3
323c09cb
602f09db
31c3200c
211c4006
32830080
12946007
32c3500c
511ca006
35830080
223c6bd2
31c30dcb
0ddb323c
3069600f
261b313c
200c600f
400631c3
0008211c
60073283
500c1494
a00632c3
0008511c
6dd23583
0ccb223c
323c31c3
600f0cdb
223c500c
323c1d0b
600f1d1b
32c3400c
31a3300c
0f8b133c
313c32c3
600f0f9b
b00c23c3
5f3225a3
0fdb323c
402c600f
1004323c
702c6ef2
0100341c
32c36ad2
602f6872
223c502c
323c1a4b
602f1a5b
313c204c
66f20014
31c3504c
081b323c
404c604f
2004323c
704c6ef2
0200341c
32c36ad2
604f6972
223c504c
323c128b
604f129b
32c3404c
31a3304c
0b0b133c
313c32c3
604f0b1b
b04c23c3
223c25a3
323c0b4b
604f0b5b
323c400c
60070404
700c1094
0040341c
32c36cd2
600f6672
20cf30cc
223c500c
323c170b
600f171b
23c370e9
0001241c
313c202c
23a30e0b
323c31c3
602f0e1b
b02c23c3
5f3225a3
0fdb323c
404c602f
304c32c3
133c31a3
32c30b8b
0b9b313c
23c3604f
25a3b04c
0bcb223c
123c13c3
204f0bdb
400631c3
000f211c
66f23283
b0ab31c3
241b353c
404c604f
304c32c3
333c31a3
233c0e4b
404f0e5b
a00632c3
0400511c
6df23583
3583704c
32c36ad2
604f7a72
223c504c
323c0ecb
604f0edb
65d2714b
23d2316b
216e614e
08040c56
40c31016
20870026
700c45b4
0d84145c
1e546007
000631c3
f000011c
40063083
3000211c
30e402c3
313c3454
6105270b
00f4233c
323c31c3
345c271b
301c0d87
311cc828
6c0c0001
0c24335c
31c303b3
211c4006
3283f000
011c0006
20c34000
175432e4
270b313c
233c60a5
31c300f4
271b323c
0d87345c
c828301c
0001311c
335c6c0c
02c30c44
36642026
00530026
08560006
00000804
0f36f016
60c3fe96
52c371c3
0d89315c
201c6732
211cc828
60070001
680c1794
21e4335c
0404435c
25a4015c
273c13c3
35c31ac0
00074664
001292dc
0d84375c
1c1b303c
0d87375c
680c0193
6de4205c
435c2037
02c30be4
404615c3
46646026
331c740b
24dc5a5a
275c0011
32c30d84
111c2006
31830007
65d2b3c3
1c0b323c
fff0b33c
c828801c
0001811c
680c28c3
6de4265c
435ce037
023c0be4
153c0020
4dc60020
46646046
640c18c3
71a4265c
435c4037
05c30e64
40062d86
466432c3
21c3376c
045402e4
740e6006
18c31bf3
435c640c
06c30c04
273c17c3
602601c0
201c4664
790022e5
25d22c09
5680763c
5840563c
c828901c
0001911c
680c29c3
0700853c
435ce037
0e060be4
201c18c3
60460120
19c34664
265c640c
403771a4
0e64435c
101c08c3
4006011c
466432c3
0c64155c
02e421c3
60060554
0046740e
355c14d3
20060484
0100111c
60073183
782c1554
0080063c
1480153c
29c36af2
335c680c
438615a4
60463664
00d3782f
680c29c3
2104335c
355c3664
341c0484
60072000
a6c35554
0c2ca21c
c828801c
0001811c
640c18c3
0984335c
17c306c3
955c3664
28c30464
e037680c
0be4435c
1ac309c3
60264046
365c4664
331c6163
0f945a5a
680c28c3
435ce037
093c0be4
301c0020
39800c2e
018e201c
46646026
c828801c
0001811c
640c18c3
71a4265c
435c4037
0ac30e64
018c101c
32c34006
365c4664
30e46dc4
28c31394
435c680c
06c320c4
2ac315c3
466437c3
68d27c0c
8580301c
2404311c
57724c0c
301c4c0f
311cc828
6c0c0001
0c04435c
17c306c3
01c0273c
46646006
22d8101c
592b7880
141c12c3
2077000f
00212f5c
78cc4c0d
0001341c
788c64d2
788f6092
08d21c0c
6672788c
11db3b3c
0006788f
786c0113
3b3c7172
786f149b
00260053
f0760296
08040f56
0736f016
90c3fe96
82c351c3
290ca3c3
1004313c
10546007
2684355c
1004233c
301c4bf2
311cc828
6c0c0001
1404335c
1a4b113c
08c33664
313c210c
60070044
355c1454
341c2684
6ff20004
c828301c
0001311c
235c6c0c
313c0a64
053c0ecb
133c0500
26640020
290c28c3
0084313c
355c6bd2
341c2684
66f20008
6186560c
4140311c
313c4c0f
6bd20104
2684355c
0010341c
562c66f2
311c6206
4c0f4140
0204313c
355c6bd2
341c2684
66f20020
6286564c
4140311c
313c4c0f
6bd20404
2684355c
0040341c
566c66f2
311c6a06
4c0f4140
341c31c3
6bd21000
2684355c
1000341c
56ec66f2
311c6006
4c0f4140
341c31c3
6bd22000
2684355c
2000341c
570c66f2
311c6086
4c0f4140
341c31c3
6bd24000
2684355c
4000341c
572c66f2
311c6706
4c0f4140
341c31c3
6ad28000
2689355c
66f26732
6786574c
4140311c
31c34c0f
411c8006
34830100
355c6dd2
34832684
301c69f2
311cc828
6c0c0001
176c6c6c
18c33664
4006650c
1000211c
68d23283
cf60201c
0001211c
6572684c
38c3684f
323c4d0c
60070804
000842dc
2681355c
60076732
32c37e94
411c8006
34830001
38546007
e007f40c
693c3594
401c5840
411cc828
700c0001
15a4335c
193c06c3
4e060500
593c3664
08c35680
29c3e00e
0f24125c
270b213c
305c09c3
323c38c4
305c271b
700c38c7
0c24335c
e08c013c
366417c3
19c3700c
38c4215c
14a4335c
e08c023c
39c33664
22e5321c
8c0d8026
68c30053
1ac0753c
32c3584c
8000341c
223c69d2
355c1c0b
323c0d84
355c1c1b
182c0d87
386c1c0f
588c3c4f
78ac5c6f
98cc7c8f
18ec9caf
790c1ccf
0003341c
301c6ed2
311cc828
6c0c0001
0d84255c
0c64335c
123c05c3
3664e08c
c828301c
0001311c
235c6c0c
355c21e4
200625a4
89ec2037
12c303c3
602627c3
00534664
790c68c3
44d22ac3
2687355c
341c0bd3
60070080
365c4254
341c0484
60070002
365c1754
760d04c1
04c9465c
065c962d
164d04d1
6272742c
301c742f
311cc828
6c0c0001
09c36eac
25c33629
742c3664
742f6172
0441165c
740c344f
0404165c
1a946027
301c34af
311c060c
6c0c4130
428b233c
0044323c
0404165c
323c6dd2
44060034
300d023c
2f5c0077
12e40021
546f0335
346f0053
0484365c
411c8006
34831000
11546007
c828301c
0001311c
265c6c0c
335c0b44
053c15a4
455c4d40
2a0025c4
36644c06
e0760296
08040f56
40c37016
d680501c
0010511c
021cc386
15c301e0
e6bc26c3
043c08cb
15c37140
e6bc26c3
0e5608cb
00000804
3f36f016
a0c3fe96
215c51c3
32c30d84
111c2006
31830800
901c63c3
65d20003
e08c623c
0001901c
56808a3c
c828701c
0001711c
b21cbac3
d01c22e6
d11c0584
c01c4130
c11c8584
355c2404
363c0d84
355c271b
340c0d87
7c0c27d2
0c24335c
200606c3
7c0c00b3
0c44335c
366406c3
0854c1a7
335c7c0c
06c30ca4
540c2026
22863664
4105111c
341c640c
60070100
2bc33594
40074809
740c3154
3cc364d2
00734c0c
440c1dc3
288c323c
00f4423c
24948027
0003341c
20546007
0424301c
4130311c
101c8c0f
111c846c
840f2404
335c7c0c
05062144
201c3664
211c0420
880f4130
8468301c
2404311c
7c0c8c0f
2144335c
00c8001c
7c0c3664
21e4235c
25a4355c
20372006
03c389ec
253c12c3
60261ac0
7c0c4664
11c4335c
15c30ac3
01c0253c
00773664
0854c1a7
335c7c0c
06c30ca4
540c2006
60573664
19946007
021c0ac3
400922e5
85c343f2
3f5c0093
600d0021
315c18c3
7b720d84
315c6f72
40260d87
040c44cf
2d540007
057302c3
335c7c0c
06c314a4
60573664
204713c3
053c0b94
101c1ac0
111cd680
43860010
08cbe6bc
921c02f3
29c3ffff
12544007
315c1ac3
931c6e04
07940001
1000341c
58c369d2
e953c1a6
0a8b333c
0010633c
0006e8b3
fc760296
08040f56
c828301c
0001311c
335c6c0c
366409c4
00000804
ff963016
105c50c3
313c6e29
203c0014
67f20340
0024313c
1d546007
5680203c
331c69cb
17945a5a
0564325c
0001341c
301c6fd2
311cc828
6c0c0001
20372006
11a4435c
123c05c3
602601c0
60264664
6e25355c
0c560196
00000804
3f36f016
70c3f796
4410c1c3
a4eca430
fff03a3c
7fa78046
0008c5dc
25c4625c
0084353c
301c6cd2
311cc828
6c0c0001
1284335c
40c33664
7b940007
67001ac3
0400933c
0024253c
51544007
821c87c3
bf3c1258
601c0140
611cc828
780c0001
15a4335c
201c0bc3
3d0022bc
36644206
101c580c
7c8022b8
425c6c0c
033c0904
208601c0
466428c3
0014353c
10546007
df5c780c
bf5c0007
40260027
8cac40b7
04000a3c
2bc319c3
466438c3
780c0153
0007bf5c
09c38ccc
28c31bc3
46643dc3
c828301c
0001311c
335c6c0c
0bc315c4
00c01c3c
36644206
0b0d303c
7f327fe5
0016233c
4f5c4137
04730081
0044353c
60078026
301c1e54
311cc828
6c0c0001
71a4175c
435c2037
09c30e64
32c31dc3
30c34664
284c2cc3
333c3103
133c0b0d
313cfff0
233cf88c
40f70016
00614f5c
099604c3
0f56fc76
00000804
3f36f016
70c3f596
040c91c3
642c00f7
a0c36137
25c4425c
6805a484
64ec6177
0204433c
c828101c
0001111c
22b8301c
80075d80
7d6c1254
0b4b033c
d7c30077
1ea0d21c
480c640c
0904335c
01c0023c
2dc32126
01d33664
d21cd7c3
640c1a88
335c480c
023c0904
210601c0
36642dc3
2ac38077
c01c682b
60270020
c01c0754
60470030
c01c0354
2dc30040
501cc8cb
511c10f8
740c0000
06c38c0c
21c32006
466431c3
740c01b7
0cc38c0c
21c32006
466431c3
801cb0c3
811cc828
48c30001
335c700c
019715a4
81572ac3
26c32a00
09c33664
341c60ec
60070010
97c37354
0e40921c
04004a3c
6f3c80b7
08c301c0
335c600c
06c315a4
22bc201c
42063d00
38c33664
721c4c0c
7c0c22b8
0904425c
01c0033c
29c32146
48c34664
401c700c
411cce0c
335c0001
04c315a4
48061ac3
08c33664
335c600c
043c1584
22060180
28c33664
c037680c
04c3accc
29c316c3
56646806
6bd26057
700c48c3
8c8cc037
02c340d7
20970805
023326c3
700c48c3
335c5c0c
023c0904
214601c0
366429c3
c037700c
00978ccc
29c316c3
46646117
c828501c
0001511c
335c740c
06c315c4
01801a3c
36644206
0007c026
740c1f94
1984435c
28060ac3
602b2bc3
740c4664
08c30193
435c600c
0ac31984
2bc32157
4664602b
680c28c3
1944435c
1cc30bc3
3dc34197
60c34664
501c6164
511c10f8
740c0000
0bc38c4c
21c32006
466431c3
8c4c740c
20060197
31c321c3
06c34664
fc760b96
08040f56
8580301c
2404311c
55724c0c
20074c0f
315c1054
341c0584
6bd20010
311c6006
215c2406
4c2f0c84
0ca4215c
01534c4f
311c6006
201c2406
211c0c00
4c2f2406
00066c4f
00000804
0336f016
91c360c3
416c82c3
2004323c
12546007
111c2006
640c4130
128b223c
308319e6
21ac323c
301c640f
311ccf30
4b260001
365c4fad
233c6e29
763c0024
a0265680
341c48f2
763c0001
52c30340
72c362f2
c828301c
0001311c
435c6c0c
06c32064
402617c3
466435c3
00470bd2
301c0994
311ccf30
0b260001
00260fcd
796c2293
211c4006
32831000
79946007
cf30301c
0001311c
0fed0b26
44d228c3
02c7383c
375c0113
173c2451
66d21f40
02c7333c
01c8321c
62863d80
4105311c
033c6c0c
00071004
984c5c94
2000441c
23948007
c828301c
0001311c
335c6c0c
06c31264
366427c3
201c0cd2
211c0604
680c4130
680f7e92
343c796c
06730f9b
0604201c
4130211c
7e72680c
796c680f
796f7e72
06d340c3
313c240c
7fa7fff0
075c25b4
640025c4
0203335c
5aa5331c
396c0554
2000141c
201c2cd2
211c0604
680c4130
680f7e72
7e72796c
0333796f
0604201c
4130211c
7e92680c
796c680f
0f9b313c
8026796f
201c01b3
211c0604
680c4130
680f7e92
303c796c
fe730f9b
501c8006
511cc828
740c0001
21a4335c
17c306c3
065c3664
30c36e29
0002341c
49546007
341c7c2c
60070004
740c1054
06c36eac
27c33e49
80273664
740c0a94
06c36eac
27c33e29
05133664
26948007
333c784c
60a7220b
301c21f4
311ccf30
4b260001
0105235c
0604201c
4130211c
7872680c
201c680f
211c8048
680c4600
680f6072
0e240116
0000041c
80560f24
00040004
14040004
001cfff3
780022da
60276c09
301c2f94
311c0608
4c0c4130
04f34e72
26948007
c800301c
0001311c
0c0f0026
2451275c
602644f2
2455375c
cf30301c
0001311c
035c0b26
301c010d
311cc828
6c0c0001
2451275c
06c38fac
60062b06
301c4664
311cc800
40060001
301c4c0f
311c8048
4c0c4600
4c0f4072
0bd209c3
c828301c
0001311c
335c6c0c
06c30fc4
00063664
0f56c076
00000804
50c33016
301c12c3
311c012c
6c0c4130
0004341c
1f546007
00a0301c
4105311c
341c6c0c
60070001
301c1654
311ccf30
4b260001
401c4ecd
411cc828
700c0001
0fe4335c
36640026
335c700c
05c30fc4
03533664
2441315c
462664f2
2445215c
cf30301c
0001311c
4eed4b26
c828301c
0001311c
215c6c0c
8fac2449
115c05c3
60062441
0c564664
00000804
40c31016
246c01c3
4e9221c3
0608301c
4130311c
31c34c0f
4000341c
201c66d2
710022da
4c0d4026
301c408c
311c060c
4c0f4130
08040856
51c37016
126412c3
25c4455c
313c4e00
758002c7
1e40433c
d00fc006
635cc88c
c84c0e47
0e67635c
635cc8ac
c86c0e87
0f47635c
640623d2
313c700f
758002c7
1e40233c
6272680c
8006680f
244d455c
655cc026
301c2455
311cc828
6c0c0001
20068e2c
31c325c3
0e564664
00000804
0336f016
80c3f896
6e29305c
09546047
0b546067
6027c006
683c0694
00730340
5680683c
00b356c3
0340683c
5680583c
18c376c3
4006656c
000f211c
80063283
0004411c
31e414c3
365c2454
341c0584
66d20001
0684265c
2627265c
301c00b3
365c5000
901c2627
911cc828
49c30001
435c700c
08c31484
400616c3
2624365c
19c34664
335c640c
08c31044
366416c3
696c28c3
0001341c
24546007
0584355c
0002341c
355c66d2
355c06a4
00f32647
5000401c
0001411c
2647455c
c828601c
0001611c
435c780c
08c31484
402615c3
2644355c
780c4664
1044335c
15c308c3
375c3664
341c0584
66d20004
06c4175c
2667175c
201c00b3
275c3000
375c2667
475c0c44
6e0025c4
1ac0873c
601cac2c
611cc828
95c30001
2000921c
275c780c
335c2664
001c15a4
011c8000
475c0001
2a0025c4
1000201c
780c3664
21e4335c
25a4275c
2026a037
80062077
8e0c80b7
13c302c3
640628c3
780c4664
21e4335c
25a4275c
101ca037
111c8000
20770001
1000401c
101c80b7
1f5c0100
80060066
20268137
81b72177
8e2c81f7
13c302c3
604628c3
375c4664
321c2664
375c1000
521c2667
59e41000
0896ba94
0f56c076
00000804
0136f016
50c3fe96
0340703c
6007626c
305c2754
341c0704
66d20040
0804205c
2787205c
600600d3
0001311c
2787305c
c828401c
0001411c
335c700c
05c31044
366417c3
2724655c
cad2c037
8e2c700c
200605c3
6f5c27c3
36c30001
653c4664
355c5680
60072c04
355c2754
341c30a4
66d20040
31a4255c
5127255c
600600d3
0001311c
5127355c
c828401c
0001411c
335c700c
05c31044
366416c3
50c4255c
4ad24077
0e30700c
200605c3
4f5c26c3
34c30021
255c8664
32c36e29
0001341c
22b8401c
63d21600
0053e00f
0296c00f
0f568076
00000804
111c2786
640c4130
e0ff201c
640f3283
22dc201c
4c0c6100
640c45d2
41ac323c
640c0093
1f00351c
6786640f
4130311c
46724c0c
08044c0f
628621c3
4105311c
341c6c0c
60070100
101c1494
111c0110
640c4130
0007241c
ff88001c
fff8011c
02c33083
323c03a3
323c202c
640f81ac
00000804
40c31016
313c01c3
60270034
66d20e54
14546047
6a946067
301c0453
311c8020
4c0c2404
00f32026
8020301c
2404311c
20464c0c
181b213c
101c0b13
111c8020
640c2404
323c4086
640f181b
0120201c
4130211c
7272680c
0913680f
8020101c
2404111c
4086640c
181b323c
201c640f
211c8014
680c2404
680f6072
22e4201c
20067100
103c2c0d
2027108b
26d21154
22542047
20942067
301c02b3
311c8620
4c0c2404
21833e06
000b251c
301c03d3
311c8624
4c0c2404
21833e06
000c251c
301c0293
311c862c
4c0c2404
21833e06
000e251c
301c0153
311c8628
4c0c2404
21833e06
000d251c
08564c0f
00000804
305c1016
67320121
62d22706
67862306
4105311c
ab10201c
0000211c
82864c0f
4105411c
23c3700c
31c32364
7bd23283
6e07205c
0121305c
43326732
323c64d2
01530034
323c2364
305c0074
60676ee7
323c0535
305c0044
08566ee7
00000804
0136f016
60c3ff96
82c351c3
400773c3
315c1754
101c2824
111cbbbb
21c30000
0a9432e4
cf30301c
0001311c
2d6d2b26
5080453c
355c03d3
65920564
315c02d3
201c26a4
211caaaa
12c30000
0a9431e4
cf30301c
0001311c
4d8d4b26
4d80453c
355c0113
64920564
0567355c
07f30026
667270ec
784c70ef
2000341c
23946007
c828301c
0001311c
335c6c0c
06c31264
25c314c3
00073664
301c1654
311ccf30
18c30001
4b2627d2
355c4dad
65920564
2b2600d3
355c2dcd
64920564
0567355c
02b30046
e0070006
301c1294
311cc828
4c0c0001
6805700c
425c6037
06c311a4
01c0153c
37c325c3
07c34664
80760196
08040f56
600764cc
315c1254
67320571
303c6ed2
113c04b0
29d23a1d
166402c3
0b0d303c
033c33c4
0053f88c
08040006
0136f016
50c3fd96
803c71c3
601c0340
611cc828
780c0001
0b24335c
780c3664
0b04435c
17c30006
30c34026
7c0c4664
000f341c
259461e7
342f2026
435c780c
01c30b04
43663c80
46646006
31c33c0c
211c4006
32830008
780c69d2
1404335c
113c05c3
40061d0b
001c3664
740022d8
21c33cab
000f241c
0f5c40b7
0c0d0041
6027742c
301c0b94
311cc828
6c0c0001
0c84335c
17c305c3
352c3664
341c31c3
60071000
313c1954
255c234b
233c0f24
5b72271b
0f27255c
000631c3
0002011c
6ad23083
148b313c
233c6025
32c31c1b
355c6f72
356c0f27
0024313c
16546007
208b313c
38c4255c
271b233c
255c5b72
313c38c7
6ad20404
11cb313c
233c6025
32c31c1b
355c6f72
d52c38c7
1000641c
1754c007
c828601c
0001611c
335c780c
05c31204
366418c3
48c3766c
4a546007
335c780c
05c30c84
366417c3
085348c3
341c756c
00260002
7a546007
5680453c
22b8101c
8c0f7480
32c3556c
011c0006
30832000
18546007
0094201c
4105211c
6172680c
401c680f
411cc828
700c0001
0fe4335c
36640026
335c700c
05c30fc4
06c33664
301c0ab3
311c012c
6c0c4130
0004341c
32c36fd2
4000341c
301c6bf2
311cc828
6c0c0001
1204335c
14c305c3
70cc3664
301c6bd2
311cc828
6c0c0001
0c84335c
17c305c3
766c3664
155c69d2
20726e29
2f5c2077
255c0021
355c6e2d
69d22c04
6e29355c
60376172
00010f5c
6e2d055c
6e29355c
600703c3
341c1954
63f20001
5680853c
c828401c
0001411c
335c700c
36642084
18c30006
98bc25c3
700c0847
1244335c
366405c3
03960006
0f568076
00000804
0336f016
50c3fd96
903c61c3
701c0340
711cc828
7c0c0001
0b24335c
7c0c3664
0b04435c
16c30006
30c34026
780c4664
000f341c
2c9461e7
342f2026
435c7c0c
01c30b04
43663880
46646006
31c3380c
211c4006
32830008
7c0c69d2
1404335c
113c05c3
40061d0b
001c3664
740022d8
21c338ab
000f241c
0f5c40b7
0c0d0041
341c788c
64d20001
6092784c
942c784f
84dc8027
301c0008
311ccf30
4b260001
301c4c0d
311cc828
6c0c0001
0c84335c
16c305c3
355c3664
341c6e04
6ef20001
0006780c
4000011c
68f23083
341c788c
04c30001
54dc6007
780c0018
0030341c
60946207
cf30301c
0001311c
4c2d4b26
c828301c
0001311c
335c6c0c
000614a4
582c3664
341c32c3
60071000
323c1a54
255c234b
233c0f24
5b72271b
0f27255c
31c3382c
011c0006
30830002
313c6ad2
6025148b
1c1b233c
6f7232c3
0f27355c
323c584c
60070024
323c1f54
255c208b
233c38c4
5b72271b
38c7255c
313c384c
6ad20404
11cb313c
233c6025
32c31c1b
355c6f72
782c38c7
1000341c
5680453c
0001801c
49c364d2
0000801c
341c782c
6bf21000
341c784c
60070002
000c62dc
49c30093
0000801c
22e6101c
4c097480
56544007
0604301c
4130311c
756f6c0c
0580301c
4130311c
752f6c0c
cf30301c
0001311c
0c4d0b26
31c3352c
1000341c
1d546007
234b313c
0f24255c
271b233c
255c5b72
31c30f27
011c0006
30830002
600749c3
313c2d54
6025148b
1c1b233c
6f7232c3
0f27355c
045349c3
303c156c
60070024
453c1d54
303c5680
255c208b
233c38c4
12c3271b
155c3b72
303c38c7
801c0404
6cd20001
11cb203c
31c34025
323c6f72
355c1c1b
801c38c7
301c0001
311cc828
6c0c0001
1204335c
14c305c3
70c33664
453c03d2
70cc5680
24546007
c828301c
0001311c
335c6c0c
05c30c84
366416c3
784cebd2
784f6172
38c4255c
270b223c
209b323c
37c3784f
600738a3
782c3c94
782f6c72
0f24255c
270b223c
235b323c
780c782f
0030341c
04546207
6192784c
784c784f
0002341c
25546007
cf30301c
0001311c
4c6d4b26
223c584c
355c208b
323c38c4
7b72271b
38c7355c
223c584c
402511cb
1c1b323c
355c6f72
301c38c7
311cc828
6c0c0001
1204335c
153c05c3
36645680
6fd2766c
cf30301c
0001311c
0c8d0b26
6e29155c
20772072
00212f5c
6e2d255c
2c04355c
301c6fd2
311ccf30
0b260001
155c0cad
21726e29
2f5c2037
255c0001
784c6e2d
0002341c
782c6bd2
1000341c
301c67f2
558022b8
5680353c
355c680f
60076e29
341c1854
63f20001
5680953c
c828401c
0001411c
335c700c
36642084
19c30006
98bc25c3
700c0847
1244335c
366405c3
6e04355c
0001341c
780c6df2
011c0006
30834000
784c67f2
0001361c
0014033c
00060053
c0760396
08040f56
2006616c
000f111c
40063183
0005211c
31e412c3
60060a94
4130311c
211c4006
4c0f0200
03f36085
211c4006
12c30004
1e9431e4
400660cc
0010211c
69d23283
311c6006
20064130
0200111c
01132c0f
311c6086
40064130
0200211c
60864c0f
4130311c
111c2006
2c0f0100
60060113
4130311c
211c4006
4c0f0300
00000804
fb96f016
d240201c
0010211c
c828301c
0001311c
68864c0f
4105311c
733c6c0c
325c094b
001c12e4
011cd800
36640001
311c6286
4c0c4105
d800301c
0001311c
6e07235c
211c4786
680c4130
0004341c
680c65f2
680f6272
301c0233
311c0580
6c0c4130
011c0006
30830800
301c67d2
311cfae6
20260001
201c2c0d
211c0094
680c4105
680f6172
311c6286
6c0c4105
0100341c
c828401c
0001411c
25546007
0604301c
4130311c
301c4c0c
311cd82c
4c0f0001
0580301c
4130311c
301c4c0c
311cd824
4c0f0001
335c700c
001c1324
011cd800
101c0001
111cd808
36640001
44dc0007
15f3003f
335c700c
001c1304
011cd800
101c0001
111cd808
36640001
08d250c3
cf30301c
0001311c
4ccd4b26
001c7bb3
011cd800
202c0001
32dc2007
301c0009
311cd80c
6c0c0001
ffff201c
07ff211c
201c3283
211cd824
680f0001
d810301c
0001311c
201c6c0c
211cffff
32830fff
d82c201c
0001211c
2027680f
700c0d94
0b04435c
101c0966
111cfae8
40460001
466435c3
205c0453
323c6e29
501c0014
511cd834
6af20001
0024323c
dd68501c
0001511c
53c363f2
afd20213
0584355c
4000341c
255c6ad2
301c0ce4
311cfae8
425c0001
8c0e025b
8580201c
2404211c
001c680c
3083f800
280c680f
d800001c
0001011c
fae8301c
0001311c
34c38c0b
07ff341c
680f31a3
6e29105c
341c31c3
6ed20001
206c612c
234b213c
323c6c72
213c235b
323c148b
7172149b
001c612f
011cd800
205c0001
32c36e29
0002341c
10546007
208c616c
208b213c
323c6172
213c209b
323c11cb
667211db
0053616f
201ca006
211cd800
686c0001
411c8006
34830100
301c6fd2
311ccf30
0b260001
684c0ced
1000101c
0001111c
727231a3
301c684f
311cfae6
4c090001
301c4bf2
311cd824
4c0c0001
0580301c
4130311c
301c0153
311c0580
4c0c4130
d824301c
0001311c
301c4c0f
311cd800
235c0001
323c6e29
66d20014
d834501c
0001511c
323c0113
65d20024
dd68501c
0001511c
355cadd2
341c0584
68d20008
d800201c
0001211c
7c72696c
401c696f
411cd800
716c0001
716f7892
301c23c3
311c0604
4c0f4130
0580201c
4130211c
7b72680c
712c680f
712f7b72
6e29345c
3e946007
cf30201c
0001211c
090d0b26
6007702c
104c2754
f004303c
13546007
220b303c
c828401c
0001411c
13d460a7
220b303c
700c60f7
1004335c
00614f5c
033304c3
341c708c
401c0001
411cc828
63d20001
0193700c
335c700c
00261004
ebf20153
c828301c
0001311c
335c6c0c
00861004
53533664
092d0b26
002652f3
24c315c3
084798bc
04dc0007
62860029
4105311c
341c6c0c
68d20100
2006706c
8000111c
60073183
301c1854
311cd800
6c6c0001
211c4006
32830100
301c6ed2
311ccf30
8b260001
6cbc8d4d
e4bc0b1b
00070b1a
0026b4dc
c828601c
0001611c
435c780c
001c2064
011cd800
15c30001
32c34006
30c34664
82dc6047
74cc0025
355c6fd2
341c0564
6ad20010
cf30301c
0001311c
2ded2b26
0624255c
401c580f
411cc828
700c0001
1444335c
d800001c
0001011c
201c3664
211cd800
682c0001
21546007
303c084c
6fd2f004
220b303c
0fd460a7
220b303c
700c6137
1004335c
00814f5c
01d304c3
341c688c
66d20001
335c700c
00861004
700c00b3
1004335c
36640026
600774cc
355c6d54
67320561
10546007
c828301c
0001311c
335c6c0c
001c15a4
011cfabc
153c0001
42060dc0
355c3664
341c0564
60071000
301c1054
311cc828
6c0c0001
15a4335c
facc001c
0001011c
0fc0153c
36644186
0564255c
8004323c
301c69d2
311cd800
055c0001
035c07c4
323c71a7
6dd20084
d800301c
0001311c
05c4155c
6e67135c
05e4455c
6ea7435c
000632c3
4000011c
69d23083
d800301c
0001311c
0604155c
6ec7135c
800632c3
0040411c
68d23483
fadc301c
0001311c
0944055c
355c0c0f
341c0584
68d20040
fae0301c
0001311c
0cc4155c
401c2c0f
411cd800
304c0001
0404313c
28546007
15c30046
98bc24c3
00070847
001954dc
341c70cc
60070020
301c1394
311ccf30
4b260001
504c4e0d
c828301c
0001311c
335c6c0c
110c19c4
170b123c
201c3664
211cd800
684c0001
684f6692
62862eb3
4105311c
341c6c0c
6cf20100
c828301c
0001311c
335c6c0c
04c313e4
260b113c
001c3664
011cd800
62290001
6fd26732
cf30301c
0001311c
8e2d8b26
c828301c
0001311c
335c6c0c
36641424
d800401c
0001411c
6e21045c
62dc0007
00660014
24c315c3
084798bc
e4dc0007
145c0013
2ad26e29
c828301c
0001311c
335c6c0c
04c31344
001c3664
011cd800
205c0001
4ad26e29
c828301c
0001311c
335c6c0c
15c313c4
62863664
4105311c
341c6c0c
60070100
101c3e54
111ccf30
6b260001
201c666d
211c0094
680c4105
680f6172
d800001c
0001011c
323c416c
60070014
32c31654
4000341c
11946007
868d8b26
c828301c
0001311c
335c6c0c
101c12c4
111cd824
25c30001
1dd33664
cf30301c
0001311c
0ead0b26
c828301c
0001311c
335c6c0c
001c1224
011cd800
36640001
15c30086
d800201c
0001211c
084798bc
24dc0007
301c000d
311c0580
6c0c4130
111c2006
31832000
1f546007
cf30301c
0001311c
4f0d4b26
0584355c
2000341c
301c6dd2
311cc828
6c0c0001
1464335c
d800001c
0001011c
301c3664
311c0580
4c0c4130
4c0f5d92
0580601c
4130611c
8006780c
4000411c
60073483
301c3054
311ccf30
0b260001
355c0f2d
341c0584
60071000
401c2454
411cc828
700c0001
001c6eac
011cd800
20060001
366425c3
335c700c
255c21e4
200625a4
80262037
20b78077
02c38e0c
253c13c3
301c1ac0
466400c7
7e92780c
0dd3780f
d800601c
0001611c
6e29065c
14540007
c828401c
0001411c
235c700c
06c30984
fab8301c
0001311c
26642c0c
335c700c
06c309e4
00a63664
201c15c3
211cd800
98bc0001
00070847
001c4994
011cd800
416c0001
0014323c
13546007
6e04305c
0001341c
241c6ed2
4bf24000
c828301c
0001311c
335c6c0c
202612a4
05d33664
15c300c6
d800201c
0001211c
084798bc
24940007
fada301c
0001311c
60276c09
301c1194
311cd800
6c4c0001
220b333c
08d460a7
0608301c
4130311c
4e724c0c
301c4c0f
311cc828
6c0c0001
1224335c
d800001c
0001011c
301c3664
311cd800
6c2c0001
e00763f2
201c1794
211cd800
682c0001
21546007
323c488c
6cd20014
800632c3
000f411c
00063483
0001011c
31e410c3
301c1294
311ccf30
4b260001
013d235c
c828301c
0001311c
335c6c0c
00260424
36642006
d800201c
0001211c
65d2682c
341c688c
69f20001
d800301c
0001311c
74a38c2c
1c94e007
cf30301c
0001311c
035c0b26
301c0145
311cc828
6c0c0001
21a4335c
d800001c
0001011c
36642006
8048201c
4600211c
6072680c
401c680f
411cc828
700c0001
1364335c
d800001c
0001011c
201c3664
211cd800
68cc0001
0020341c
15946007
313c284c
60070404
301c1054
311ccf30
0b260001
014d035c
335c700c
090c19c4
170b113c
01f33664
fada301c
0001311c
60276c09
301c0894
311c0608
4c0c4130
4c0f4e72
c828301c
0001311c
335c6c0c
001c07a4
011cd800
36640001
0f560596
00000804
fa967016
21772006
00404f3c
01405f3c
403740c6
101c04c3
111cc800
301c0001
311cd5e8
4ca00001
1abc35c3
60c60878
04c36037
d800101c
0001111c
22ec201c
1abc35c3
001c0878
011cc000
101c0001
111c0120
301c0010
311cc130
4c200001
08cbb0bc
24060006
0010111c
0100201c
08cbb0bc
13a0001c
0000011c
1478301c
0000311c
9cbc2c20
48bc08cb
301c0860
311ccf30
233c0001
89c602f0
00df433c
fc9432e4
2c0d2006
084b06bc
06960006
08040e56
40c33016
0094301c
4040311c
341c6c0b
6df20001
c828301c
0001311c
335c6c0c
00062164
9000011c
36643fe6
80bc0006
82200895
c828501c
0001511c
00040004
00040004
335c740c
00062184
62203664
f5d46007
08040c56
40c33016
21af2006
211c4006
205c0400
60062767
1000311c
2747305c
620f6406
4006624f
0001211c
2787205c
105c2026
20062b47
0800111c
5107105c
111c2006
105c1200
305c50e7
205c2ba7
301c5127
418022b8
0340303c
101c680f
111caae5
105cd95e
301c71a7
311c4800
305c01e8
201c6e67
211cb400
205c04c4
305c6e87
301c6ea7
305c733c
101c6ec7
008022bc
42062686
0891b0bc
22cc201c
21861100
b0bc4186
501c0891
511cc828
740c0001
045c6c6c
36646e84
335c740c
04c311e4
740c3664
d69c101c
0010111c
21e7135c
08040c56
226420c3
0610001c
4130011c
6026200c
31a33223
0804600f
326430c3
1000201c
1180211c
233c6d00
680c100c
680f6772
6692680c
0804680f
326430c3
1000201c
1180211c
233c6d00
680c100c
680f6472
00000804
211c4006
680c4130
0804680f
326430c3
1000201c
1180211c
233c6d00
680c100c
ff3f341c
31ac313c
680f3364
00000804
326430c3
1000201c
1180211c
233c6d00
680c100c
fffc341c
336431a3
0804680f
326430c3
100c213c
1000101c
1180111c
133c6c80
640c100c
fffb341c
03fc241c
640f32a3
00000804
326430c3
180c213c
1000101c
1180111c
133c6c80
640c100c
fff7341c
07f8241c
640f32a3
00000804
326430c3
200c213c
1000101c
1180111c
133c6c80
640c100c
ffef341c
0ff0241c
640f32a3
00000804
326430c3
280c213c
1000101c
1180111c
133c6c80
640c100c
ffdf341c
1fe0241c
640f32a3
00000804
311c6006
201c4140
4c0f2000
40066705
1000211c
08044c0f
311c6006
201c4140
4c0f4000
00000804
311c6006
201c4140
211c2000
4c0f0002
00000804
400f4026
00000804
03c3604c
00000804
606f642c
00000804
40af43e6
241c444c
408f001f
00000804
40ef4026
40cf446c
40ef4046
00000804
65d264cc
610f6086
007360ef
610f6086
00000804
341c648c
60270007
60470954
60071054
64061894
4806616f
640602f3
4806614f
648c416f
28cb333c
01f3614f
616f6406
414f4806
333c648c
7fe5220b
00b3618f
616f6806
416f4406
00000804
311c6006
616fff00
64326629
614f7812
7c12652b
0804614f
341c648c
60470007
604c0594
0002341c
604c7dd2
0001341c
61cc7dd2
400f4026
080403c3
401c3016
411ccf60
704c0001
323c43e6
704f281b
6006102f
708c706f
182b333c
00f8351c
323c4086
4046221b
231b323c
323c4106
708f241b
70ef6006
6026710f
600670cf
501c716f
511cc828
740c0001
0d04335c
740c3664
0d64335c
0800001c
2040011c
366414c3
335c740c
001c0d84
011c0800
14c32040
740c3664
0da4335c
0800001c
2040011c
366414c3
335c740c
001c0dc4
011c0800
14c32040
740c3664
0de4335c
0800001c
2040011c
366414c3
335c740c
001c0e04
011c0800
14c32040
201c3664
211c0800
301c2040
696f0080
64d270ec
0080301c
0c56694f
00000804
0136f016
60c3fb96
72c341c3
02d753c3
cf60301c
0001311c
21c32c2c
095402e4
c828301c
0001311c
335c6c0c
36640e44
0030243c
23837f86
0030453c
101c4383
111ccf60
644c0001
0020341c
1c546007
20c64cd2
0f3c2037
16c30040
0824301c
2040311c
085d72bc
46548007
403740c6
00400f3c
24c317c3
0824301c
2040311c
085d72bc
052b0733
341c30c3
533c000f
86c3100c
0800601c
2040611c
12c30273
023525e4
79ac15c3
0004341c
31c37df2
08c300f3
0004821c
192f000c
7af27f85
400748a0
17c3ed94
0800201c
2040211c
04c30233
023545e4
69ac05c3
0004341c
30c37df2
613c00b3
c92f024f
7cf27f85
80079020
301cef94
311cc828
6c0c0001
0e24335c
0800001c
2040011c
cf60101c
0001111c
05963664
0f568076
00000804
22642412
0ff0141c
44124880
440c2100
209b233c
0804440f
0736f016
90c3ff96
00d7313c
c018001c
0001011c
101cac00
111cc04c
ec800001
c080201c
0001211c
8006cd00
c828a01c
0001a11c
0b1385c3
60377809
00ff331c
1ac30954
335c640c
2f5c0e84
02c30001
343c3664
6087ffc0
80a735b4
28c31b94
04092a00
1000201c
1180211c
233c6100
680c100c
ff3f001c
680f3083
001c4409
011c1000
68001180
100c233c
6672680c
34090313
1000201c
1180211c
233c6500
680c100c
ff3f001c
680f3083
201c3409
211c1000
65001180
100c233c
6772680c
0006680f
4613011c
54092006
009f373c
085328bc
600c0ac3
0ea4335c
009f053c
80253664
61a6c025
22f219c3
43e46126
0196a474
0f56e076
00000804
211c4006
680c4600
111c2006
31a30700
4205680f
7a72680c
0804680f
211c4086
680c4600
111c2006
31a30700
0804680f
40c31016
0200041c
085334bc
0853b2bc
311c6006
8c0f4617
08560006
00000804
0736f016
80c3fc96
a2c391c3
0080433c
f06bd04b
c828501c
0001511c
335c740c
36640ce4
343c540c
60370080
00266f5c
0080363c
60b77180
00667f5c
1964425c
19c308c3
36c32ac3
04964664
0f56e076
00000804
fc96f016
01436f5c
01835f5c
c828401c
0001411c
e2d7900c
5f5ce037
00b70026
00661f5c
19a4445c
13c302c3
36c34257
04964664
08040f56
0336f016
81c370c3
336492c3
2a546047
4f546067
7d946027
10f8601c
0000611c
8c0c780c
20060d86
31c321c3
50c34664
c828401c
0001411c
335c700c
2d861584
700c3664
1764335c
366405c3
335c700c
05c31784
28c317c3
700c3664
17a4335c
601c09d3
611c10f8
780c0000
001c8c0c
200600cc
31c321c3
50c34664
c828401c
0001411c
335c700c
101c1584
366400cc
335c700c
05c317c4
700c3664
17e4335c
17c305c3
366428c3
335c700c
04f31804
10f8601c
0000611c
8c0c780c
00cc001c
21c32006
466431c3
401c50c3
411cc828
700c0001
1584335c
00cc101c
700c3664
1824335c
366405c3
335c700c
05c31844
28c317c3
700c3664
1864335c
19c305c3
780c3664
05c38c4c
21c32006
466431c3
c0760006
08040f56
3f36f016
d0c3a696
c2c32077
0ce4bf5c
936493c3
0cc3af5c
0d037f5c
c828501c
0001511c
8f3c740c
335c1040
08c31584
36642c86
335c740c
0f3c1584
2c860a00
740c3664
00806f3c
1584335c
101c06c3
36640098
335c740c
06c31724
36642006
ff47301c
54940007
c037740c
1744435c
19c30cc3
3ac35957
00074664
e8073f94
740c0894
1884435c
18c4335c
02530086
0894e407
435c740c
335c1884
004618c4
e6070133
740c2b94
1884435c
18c4335c
366400a6
08c330c3
27c31bc3
50c34664
c828701c
0001711c
8f3c7c0c
6f3c0a00
c0370080
18a4435c
20570dc3
6c8628c3
05e44664
7c0c0b94
15c4335c
1f3c08c3
25c31040
40c33664
06c307d2
0b1ce6bc
ff47301c
06c300b3
0b1ce6bc
03c334c3
fc765a96
08040f56
301c3016
311c0608
6c0c4130
0400341c
ff35001c
34946007
301c03c3
311cd800
135c0001
200771c1
301c2b94
311cfab8
4c0c0001
0564325c
0400341c
2000501c
525c63d2
401c07a4
411cc828
700c0001
0cc4335c
301c3664
311cfab8
4c0c0001
335c700c
125c1664
148025c4
301c3664
311cd800
40260001
71c5235c
0c560006
00000804
41c31016
0b64205c
1b544007
fab8301c
0001311c
305c0c0c
298025c4
331c640b
0f945658
32c3442b
341c3443
69d20001
0010343c
3a1d313c
25c4205c
00530d00
08560006
00000804
0736f016
fba8f21c
31c380c3
326462c3
0f3c62b7
20064440
bebc4206
1fe60891
200718c3
001bf2dc
01413f5c
901c3064
39e40000
62970815
041c03c3
02b7007f
0080901c
22977809
32e421c3
18290894
341c30c3
60070002
0019c4dc
c828401c
0001411c
335c700c
08c308e4
36642297
1fc670c3
62dce007
700c0019
1584335c
02c00f3c
0418101c
22973664
5fe521c3
3f5c4277
60270121
22970835
410721c3
01c30454
50940127
21c32297
06944027
60277c09
001704dc
22970373
410721c3
7c090694
74dc6107
02530016
21c32297
06944047
60477c09
0015e4dc
22970133
412721c3
7c090594
54dc6127
3c290015
0014313c
e2dc6007
501c000a
511cc828
740c0001
188c013c
435c0237
08c30924
01012f5c
400612c3
45403f3c
30c34664
b3dc6007
20260013
016d1f5c
22a32f5c
01762f5c
1c2b740c
20060037
20b72077
01c38cec
22971013
40a721c3
0011f2dc
31c301c3
000a361c
133c7fe5
30c3f88c
61f77fa5
00e13f5c
04356027
12dc2007
5c09000e
06544067
30c30297
b2dc6067
41470010
20070454
001064dc
31c32297
0004361c
7f327fe5
04544087
b4dc6007
3c29000f
0044513c
2354a007
60071f26
000f92dc
42725829
3f5c41b7
782d00c1
c828301c
0001311c
213c6c0c
4177188c
0924435c
3f5c08c3
13c300a1
417229c3
45403f3c
30c34664
38dc6007
1ab3000d
0014313c
2e546007
c828901c
0001911c
680c29c3
188c213c
435c4137
08c30924
00813f5c
25c313c3
45403f3c
30c34664
b3dc6007
2026000b
016d1f5c
22a32f5c
01762f5c
600c09c3
20373c2b
a0b7a077
05c38cec
0180173c
0080263c
02c03f3c
313c04d3
401c0024
411cc828
60070001
301c2054
311cfab8
4c0c0001
5f3c700c
335c02c0
023c0904
20c601c0
366425c3
d4dc0007
700c0008
20373c2b
00b70077
173c8cec
263c0180
35c30080
01534664
335c700c
063c15a4
173c0080
5c2b0180
901c3664
911cc828
29c30001
af3c680c
335c02c0
0ac31584
0418101c
301c3664
311cfab8
4c0c0001
600c09c3
0904335c
01c0023c
2ac320c6
00073664
19c35894
875c640c
5f3c0013
a0374440
063c8ccc
101c0080
111cfabc
2ac30001
466438c3
680c29c3
15c4335c
173c05c3
42060080
00073664
7c2b3e94
1c2c782e
05d3182f
21c32297
2a9440c7
60c77c09
3c292c94
0044313c
15546007
013c700c
00f7188c
0924435c
2f5c08c3
12c30061
3f3c4006
46644540
600730c3
20261874
0153382d
335c700c
063c15a4
173c0080
5c2b0180
5c2b3664
7c2c582e
0f5c782f
180d0141
01130006
00d31fa6
00931f86
00531f66
f21c1f46
e0760458
08040f56
ff96f016
73c34037
626461c3
c828501c
0001511c
335c740c
20a608e4
40c33664
80071fe6
740c1c54
1644335c
30c33664
60071f26
540c1474
0040143c
02c7363c
16c4425c
20060580
00013f5c
37c323c3
30c34664
60071f46
00060274
0f560196
00000804
3f36f016
f398f21c
c1c390c3
0fc362c3
0c54021c
42062006
0891bebc
43375889
01c07c3c
501ce2f7
511cc828
740c0001
08e4335c
12c307c3
b0c33664
1bc31fe6
12dc2007
740c0031
1584335c
46400f3c
0418101c
740c3664
15a4335c
021c0fc3
19c30c54
22bc121c
36644206
30c30317
60277fe5
000ce5dc
335c740c
0f3c1584
101c03c0
36640428
2bc3784c
07c3e82c
c9dc30e4
2317002d
402721c3
3f5c0694
3f5c0181
009301e5
7f5ce046
801c01e5
811cc828
08c30001
39c3400c
22b8321c
df3c6c0c
425c4640
033c0904
20c601c0
46642dc3
000770c3
002bb4dc
01c0a63c
4c0c38c3
3fc3b86b
0c54321c
88cc6037
19c30ac3
22bc121c
35c32dc3
08c34664
335c600c
0f3c15a4
1fc30440
0c54121c
36644206
513c38a9
abd20024
600c08c3
2037386b
4026e077
8cec40b7
053307c3
0014313c
2b546007
7c0c78c3
188c213c
435c4277
02d70924
01213f5c
25c313c3
321c3fc3
46640c64
600730c3
0027b3dc
1f5c2026
2f5c232d
2f5c6323
78c32336
186b7c0c
a0770037
20b72026
05c38cec
2f3c1ac3
3dc30540
01f34664
0044313c
24dc6007
28c30026
335c680c
0f3c15a4
1ac30540
3664586b
3f5c7889
f8a901e5
01ed7f5c
0f5c186b
384c01f6
501c2437
511cc828
740c0001
0428201c
701c4037
e0775aa5
0964435c
1cc309c3
3f3c2bc3
466403c0
000740c3
002314dc
10c30317
08942027
335c740c
09c31584
1a88021c
740c4413
1584335c
021c09c3
43331ea0
10c30317
559420a7
433258a9
1f4643b7
15dc4267
740c0022
a21cafc3
335c087c
0ac31584
0374101c
0f5c3664
0f5c0181
8fc343e5
0880821c
335c740c
08c315a4
00401b3c
0370201c
740c3664
1644335c
00073664
001fb3dc
7fc3740c
0c28721c
1684435c
01c0063c
01c12f5c
586b12c3
37c34312
30c34664
a3dc6007
740c001e
213c2397
335c02c7
18c315a4
17c30500
36644586
201c740c
40370374
5aa5701c
435ce077
09c30964
2bc31cc3
11533ac3
30c30317
0007361c
233c7fe5
42b7f88c
7fa530c3
04356027
f2dc4007
301c0014
311cc828
6c0c0001
1584335c
03c00f3c
0428101c
23173664
406721c3
784c0894
1c2c7bc3
31e410c3
001a19dc
733c78a9
e377188c
0004341c
61546007
30c30317
0004361c
533c7fe5
a5f2f88c
20072297
001932dc
43124357
3f5c4237
78ad0101
f88de0a6
c828401c
0001411c
335c700c
09c30944
26c31cc3
00073664
001814dc
6f3c700c
335c03c0
0f3c1584
101c0540
36640410
02720217
1f5c01f7
1f5c00e1
458601ed
01f62f5c
1054a007
3f5c6086
700c01e5
e037e706
5aa5001c
435c0077
09c30964
2bc31cc3
20e60293
01e51f5c
e357700c
4287273c
0428001c
101c0037
20775aa5
0964435c
1cc309c3
4d003bc3
466436c3
a4dc0007
28930013
c828801c
0001811c
5c0c78c3
321c39c3
6c0c22b8
4640df3c
0904425c
01c0033c
2dc320c6
70c34664
44dc0007
a63c0012
18c301c0
b86b440c
321c3fc3
60370c54
0ac388cc
121c19c3
2dc322bc
466435c3
600c08c3
15a4335c
04400f3c
121c1fc3
42060c54
38a93664
0024513c
08c3abd2
386b600c
e0772037
40b74026
07c38cec
313c0533
60070014
78c32b54
213c7c0c
41b7188c
0924435c
3f5c02d7
13c300c1
3fc325c3
0c64321c
30c34664
43dc6007
2026000e
232d1f5c
63232f5c
23362f5c
7c0c78c3
0037186b
2026a077
8cec20b7
1ac305c3
05402f3c
46643dc3
28c30153
335c680c
0f3c15a4
1ac30540
3664586b
3f5c7889
f8a901e5
01ed7f5c
0f5c186b
384c01f6
501c2437
511cc828
6f3c0001
429703c0
16544007
e357740c
4287273c
0428001c
101c0037
20775aa5
0964435c
1cc309c3
4d003bc3
466436c3
21540007
740c12f3
e037e706
5aa5001c
435c0077
09c30964
2bc31cc3
466436c3
84dc0007
23170008
406721c3
740c0c94
1584335c
021c09c3
101c0e40
36640418
10b30297
c828301c
0001311c
335c6c0c
09c31584
1258021c
0418101c
0ed33664
32c34317
6e9460c7
335c740c
0fc31584
0bf0021c
36642706
133c78a9
21770044
24542007
0f84733c
0f5ce137
18ad0081
388d20a6
335c740c
09c30944
26c31cc3
00073664
740c5194
1584335c
021c0fc3
24060c08
65863664
5f963f5c
e0f7e272
00617f5c
5f8d7f5c
740c0253
15a4335c
021c0fc3
163c0c08
586b01c0
586b3664
5f962f5c
00a13f5c
5f8d3f5c
321c3fc3
00c60c68
c45e033c
c828501c
0001511c
2706540c
701c2037
e0775aa5
0964425c
1cc309c3
46642bc3
0cf240c3
335c740c
09c31584
1670021c
0418101c
04c33664
1ee601d3
1fc60193
1fa60153
1f860113
1f0600d3
1f260093
00060053
0c68f21c
0f56fc76
00000804
fe963016
215c52c3
60260544
14544007
c828301c
0001311c
401c6c0c
80370190
4aa4401c
435c8077
353c0964
466401c0
02f27ee6
03c330c3
0c560296
00000804
0f36f016
b0c3f896
42c351c3
642c63c3
0004341c
301c6ad2
311cc828
6c0c0001
26096eac
366425c3
8000a01c
0001a11c
1ac34497
7fe7215c
301c84c3
8383f000
7fc7815c
c828901c
0001911c
640c19c3
15a4335c
18c30ac3
0ff8201c
29c33664
243c680c
335cfff4
1ac315a4
16c30880
36644457
680c29c3
21e4235c
1ac0753c
25a4155c
7112746c
d000321c
60266037
60066077
8a0c60b7
12c301c3
640627c3
19c34664
235c640c
155c21e4
746c25a4
321c7112
6037d000
0027af5c
1000301c
301c60b7
3f5c0100
60060066
60266137
60066177
602661b7
8a2c61f7
12c301c3
604627c3
60c34664
53940007
640c19c3
21e4335c
25a4255c
00078f5c
20772026
8e0c00b7
13c302c3
640627c3
29c34664
335c680c
255c21e4
8f5c25a4
af5c0007
101c0027
20b71000
0100101c
00661f5c
2026c137
c1b72177
8e2c21f7
13c302c3
604627c3
60c34664
23940007
680c29c3
21e4235c
25a4155c
7112746c
d000321c
60266037
00b76077
01c38a0c
27c312c3
46646406
341c742c
03c30004
19c36bd2
6eac640c
36290bc3
366425c3
005306c3
08960026
0f56f076
00000804
1f36f016
90c3f896
a03c61c3
c01c5680
c11ccf30
801c0001
811cc828
b01c0001
b11c8000
165c0001
786c25c4
6c807112
dffc321c
32c34c0c
ccaa361c
0b0d333c
7f327fe5
5aa5231c
64f20554
4aa4231c
0b267a94
0b4d2cc3
12546007
0564365c
211c4006
32831000
f000701c
0000711c
765c6dd2
301c0c24
7383f000
786c00f3
6c807112
dff8321c
08c3ec0c
121c400c
786cd000
425c7112
001c15a4
011c8000
25800001
0ff8201c
40064664
215c1bc3
215c7fc7
08c37fe7
235c600c
563c21e4
365c1ac0
e03725a4
20772026
00b70006
03c38a0c
25c312c3
46646406
640c18c3
21e4335c
25a4265c
001ce037
011c8000
00770001
1000101c
001c20b7
0f5c0100
20060066
00262137
21b70177
8e2c21f7
13c302c3
604625c3
18c34664
235c640c
165c21e4
786c25a4
321c7112
6037d000
60776026
00b70006
01c38a0c
25c312c3
46646406
215c19c3
32c36e29
0003341c
06946067
6027780c
6ac30354
0896ecb3
0f56f876
00000804
6ee4305c
0e946047
cf94301c
0001311c
0200233c
23c34cef
0380101c
a020111c
602701f3
301c1194
311ccf94
233c0001
4cef0200
101c23c3
111c0080
123ca020
4c6f087e
101c2c0f
111ccf94
21c30001
301c2364
311c0080
4c0e2100
808c213c
4c0e6045
00000804
40c33016
215c01c3
40476ee4
01731894
341c680c
6dd2a000
341c680c
68a700ff
08b30894
111c2346
46862020
4105211c
341c640b
60070004
03f3ec94
40272006
60862894
2020311c
61054c0e
20064c0e
2020111c
211c4686
01534105
341c680c
66d2a000
341c680c
68a700ff
640b2054
0001341c
00f374d2
0380301c
2020311c
00f32c0c
311c6306
6c0b2020
136413c3
c828301c
0001311c
335c6c0c
24c30844
60063664
2020311c
4c0e4026
08040c56
c0963016
205c52c3
40476ee4
141c0994
013c1fff
3f860030
80260183
800601b3
402704c3
141c0994
013c1fff
101c0ff0
0183ff00
323c42c3
6027fff0
301c2bb4
311ccf94
a7d20001
101cec31
111c9000
00d30001
101cec31
111c8000
2caf0001
06944047
e80c343c
00c5233c
402700f3
343c0a94
23c3e80c
301c4872
311ccf94
4c4f0001
e82c243c
cf94301c
0001311c
201c4ccf
211ccf94
68cc0001
68cf6e72
311c6146
201c2100
4c0e0085
211c41c6
680b2100
0004341c
61c67dd2
2100311c
2c0e2086
0c564096
00000804
0336f016
90c3fe96
61c383c3
0030423c
42835f86
733c6257
0373c005
431c54c3
03351f00
1f00501c
0081201c
35c34037
1fff341c
4000201c
1488211c
607732a3
17c309c3
38c326c3
08772abc
da8092a0
e5948007
c0760296
08040f56
22642412
0ff0141c
44124880
440c2100
209b233c
0804440f
0136f016
70c3fd96
62c351c3
8f5c23c3
301c0124
311cc828
6c0c0001
21e4135c
38c3854c
25a4035c
02944047
a0374066
c0b74077
1ac0283c
466437c3
80760396
08040f56
31c31016
326412c3
00474606
00471054
406607b4
41260cd2
08940027
46e60113
05540067
008747a6
40060254
13542007
1000101c
1180111c
67d24880
680c4212
ff3f401c
02333483
680c4212
ff3f101c
02933183
411c8006
4a00104e
42126ad2
101c680c
3183ff3f
680c680f
00d36772
680c4212
ff3f401c
680f3483
08040856
004745c6
00470e54
40c605b4
08940027
46860113
05540067
00874746
40060254
011c0006
6800104e
100c133c
011c0006
68002010
080c033c
640c4006
313c6492
6406027f
016f303c
40c74025
0804f794
0087f016
00871e54
45c60fb4
8026a006
004765c3
46864a54
47b40047
806640c6
3e940027
00c70853
40061154
8026a746
00c7c046
00e73a14
01a70e54
01b33194
a0064746
65c38046
20c30613
8066a746
0573c046
053345c6
81b4301c
4600311c
301c8c0f
311c6000
4c0f4600
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
2198321c
ec0fe106
000606f3
50c320c3
60c38026
16942007
711ce006
6b802010
080c733c
311c6006
4980104e
43644212
016f473c
6472680c
027f323c
20c72025
0087f894
40061935
2010211c
433c7500
e006080c
104e711c
133c7780
4006100c
036406c3
016f043c
6472640c
027f313c
40c74025
0f56f894
00000804
f8967016
51c300f7
211c4106
680c4600
1800351c
20c3680f
608730c3
60c36d54
0db44087
3054c027
000720c3
40472054
20c33f54
a4dc4067
0993000f
63c360d7
b2dcc147
23c30009
08b46147
410762c3
c1276054
000eb4dc
40d70e73
618732c3
000a82dc
24dc41a7
1773000e
c828301c
0001311c
335c6c0c
6f5c0e84
06c30061
40d73664
401c1bd3
411cc828
700c0001
0e84335c
00616f5c
366406c3
335c700c
00460e84
40c63664
61464137
401c1993
411cc828
700c0001
0e84335c
36640166
335c700c
01860e84
c5c63664
4146c137
401c10d3
411cc828
700c0001
0e84335c
366401a6
335c700c
01c60e84
66863664
c0466137
301c0813
311cc828
6c0c0001
0e84335c
366401e6
41374746
13736046
c828401c
0001411c
335c700c
00060e84
700c3664
0e84335c
366401a6
335c700c
01c60e84
c0063664
4026c137
401c0a13
411cc828
700c0001
0e84335c
36640026
335c700c
00460e84
700c3664
0e84335c
366401a6
335c700c
01c60e84
60c63664
c1466137
0d13c177
c828401c
0001411c
335c700c
01660e84
700c3664
0e84335c
36640186
335c700c
01a60e84
700c3664
0e84335c
366401c6
413745c6
097360d7
c828401c
0001411c
335c700c
01e60e84
700c3664
0e84335c
366401a6
335c700c
01c60e84
c7463664
4046c137
06934177
81b4301c
4600311c
cc0fc026
6000301c
4600311c
4c0f4006
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
4c0f6085
2198321c
cc0fc106
301c0b93
311cc828
6c0c0001
0e84335c
36640006
40f74006
60264137
a0076177
6f5c2894
c1f70081
c828501c
0001511c
c037c0c5
00014f5c
011c0006
20064613
00e13f5c
6f5c23c3
36c300a1
085da0bc
335c740c
2f5c0ea4
02c300e1
61d73664
c02563c3
2f5cc0b7
41f70041
e59424e4
26c3c0d7
21354087
61b76686
c828401c
0001411c
011c0006
20064613
00c16f5c
614626c3
085da0bc
335c700c
2f5c0ea4
02c300c1
61973664
c02563c3
2f5cc077
41b70021
e7944747
0e560896
00000804
0580301c
4130311c
02c34c69
0001041c
00000804
0860ccbc
00000804
0860c4bc
00000804
0860d4bc
00000804
086060bc
d024301c
0001311c
5800201c
0001211c
001c4c0f
b6bc2800
08040860
cf30301c
0001311c
235c4b26
08040165
301c1016
311c10f8
101c0000
111c7d1c
2c0f0016
10fc401c
0000411c
cfb4301c
0001311c
03c3700f
9cbc2e06
700c08cb
4c0f4006
2c8d2006
4cad4026
41064ccd
4d0d4ced
4d2d40c6
1478201c
0000211c
280f2006
c0b0201c
0010211c
4c8f4c6f
101c4caf
111cc064
2ccf0010
4d0f4cef
4d4f4d2f
c164101c
0010111c
4d8f2d6f
4dcf4daf
4e0f4def
4e4f4e2f
4e8f4e6f
4ecf4eaf
4f0f4eef
4f4f4f2f
08564f6f
00000804
001302f2
00000804
301c20c3
311cd024
6c0c0001
03c36065
01833f86
2cbc12c3
08040a80
0a80c4bc
00000804
0860c4bc
00000804
5cbc03d2
08040a7f
0860ccbc
00000804
0a7e8abc
00000804
0860d4bc
00000804
08040013
00000804
00000804
00000804
00000804
0b64105c
301c640f
6d200200
644e3364
646e6026
23c364eb
48f22364
644f640c
3364644b
444e64ee
0804446e
00000804
d02c301c
0001311c
4c0f4006
00000804
305c6046
080405ed
fc963016
01002f3c
ffde023c
0b00301c
501c0c0c
511cd02c
60260001
301c740f
311cc828
2c0c0001
311c6006
60370002
0e64305c
00c0321c
60266077
00463f5c
1e24415c
402612c3
46646066
7ff2740c
0c560496
00000804
0b00301c
6abc0c0c
080408bb
fd967016
40e750c3
201c3394
211cd030
301c0001
311cd038
680f0001
d238101c
0001111c
305c282f
60a70b89
305c2194
6c8c0b24
1c946007
62c343c3
363c02b3
40464a1d
255c4037
221c0e64
40770080
1f5c2026
05c30046
201c13c3
60460200
08d1babc
355c8025
43e405e9
0396e974
08040e56
fd963016
341c612c
60070001
301c2254
311ccf30
4b260001
015d235c
0e00501c
4130511c
433c740c
940f0115
233c612c
2264164b
033c4037
133c084b
233c088b
333c08cb
74bc190b
7dc6088f
940f4383
0c560396
00000804
60c37016
d800301c
0001311c
6e29235c
0014323c
d834501c
0001511c
323c6af2
60070024
000c72dc
dd68501c
0001511c
d800301c
0001311c
6ee4335c
608754cc
4fd22094
0569355c
6bd26732
0f80463c
155c04c3
42460884
08cbb0bc
08c7465c
600774cc
355c3654
40060564
0001211c
60073283
463c2e54
355c1200
045308a4
12544007
0564355c
111c2006
31830002
463c6bd2
04c30f80
08c4155c
b0bc4246
465c08cb
74cc08c7
13546007
0564355c
211c4006
32830004
463c6cd2
355c1200
04c308e4
4c2b13c3
08cbb0bc
08e7465c
d800201c
0001211c
6007682c
69cb1a54
17546007
200729eb
463c1454
04c30f80
08c4165c
b0bc4246
063c08cb
101c1000
111cd81c
40860001
08cbb0bc
08c7465c
600774cc
355c1854
40060564
0008211c
60073283
001c1054
011cd58c
155c0001
41460904
08cbb0bc
d58c301c
0001311c
0867365c
600774cc
355c1854
20060564
0010111c
60073183
001c1054
011cd598
155c0001
47860924
08cbb0bc
d598201c
0001211c
0887265c
d800201c
0001211c
6007682c
686c1754
111c2006
31830800
06c364d2
08be46bc
d800301c
0001311c
40066c6c
1000211c
64d23283
d8bc06c3
0e5608bc
00000804
ff961016
305c40c3
63270649
000b64dc
0653305c
72546667
07b46667
0f546227
f4dc6447
0713000a
22dc6aa7
6cc70008
0008c2dc
54dc6887
0db3000a
12dc2007
305c000a
60870673
0009c5dc
08946087
311c6786
2c0c4105
0547105c
604701d3
67860694
4105311c
00b36c0b
311c6786
6c094105
0547345c
200604c3
0a80243c
0673345c
08bc6cbc
200604c3
32c34006
08bb50bc
20070ed3
66861454
4105311c
0567305c
105c2006
305c05a7
60870673
202668b4
05a7105c
203c2006
0a930b00
05a4305c
5d546007
05a7105c
0673305c
07946087
0564305c
0584105c
0a332c0f
0564205c
0584405c
60478037
880e0394
3f5c0913
680d0001
20070893
305c4254
331c0673
3db41000
201c2006
211c8000
05530001
35542007
0673305c
1000331c
200630b4
9000201c
0001211c
200703b3
205c2854
231c0663
23b40fff
301c2006
311c8000
01b30001
1b542007
0663205c
0fff231c
200616b4
9000301c
0001311c
345c4980
50bc0673
04c308bb
40062006
6cbc32c3
00b308bc
21c32006
08b7e2bc
08560196
00000804
fe96f016
61c370c3
a0466364
00055f5c
4f5c8026
20860025
600626c3
08bbcabc
00055f5c
00254f5c
208607c3
34c326c3
08bbcabc
00055f5c
00254f5c
20a607c3
600626c3
08bbcabc
00055f5c
00254f5c
20a607c3
34c326c3
08bbcabc
0f560296
00000804
60c37016
6e29105c
341c31c3
203c0001
63d25680
0340203c
6bd268cc
0564325c
4000341c
425c66d2
525c0844
01330864
bc00401c
0001411c
0800501c
0000511c
d028301c
0001311c
4c0d4026
0b00301c
04c38c0f
01d4101c
08cb9cbc
0e67545c
3000353c
0e87345c
0e47445c
1d40343c
0e27345c
6ee1365c
0b8d345c
145c2006
001c0b85
011cd4f8
2d860001
08cb9cbc
d4f8201c
0001211c
0b27245c
c0d8301c
0001311c
0b47345c
145c2006
404605c7
05ed245c
0b89345c
079460a7
d564201c
0001211c
0b67245c
d438001c
0001011c
00c0101c
08cb9cbc
d4f8301c
0001311c
d438101c
0001111c
345c2c0f
44060b24
101c4ece
111c0800
2caf0002
c0b4201c
0001211c
0e07245c
0b89345c
069460a7
cb64301c
0011311c
301c684f
311cd4f8
2c0c0001
0200313c
4c2f4046
245c4c4f
221c0e64
4c6f0080
4c8f4066
211c4006
4caf0002
0e64245c
00c0221c
40064ccf
4dee4dce
0400313c
4c2f4086
245c4c4f
221c0e64
4c6f0100
4c8f40a6
211c4006
4caf0004
0e64245c
0140221c
40064ccf
40464dce
313c4dee
40c60600
41064c2f
245c4c4f
221c0e64
4c6f0180
4c8f40e6
211c4006
4caf0008
0e64245c
01c0221c
40064ccf
4dee4dce
0800313c
4c2f4106
4c4f4206
0e64245c
0200221c
41264c6f
40064c8f
0010211c
245c4caf
221c0e64
4ccf0240
4dce4006
313c4dee
21460a00
44062c2f
245c4c4f
221c0e64
4c6f0280
2c8f2166
211c4006
4caf0020
0e64245c
02c0221c
20064ccf
2dee2dce
08040e56
65530a0d
5220646e
31313953
424e2e36
43572e5a
4e45472e
2e782e52
2e782e78
0d737072
0000000a
65530a0d
5220646e
31313953
424e2e36
344d2e5a
4e45472e
2e782e52
2e782e78
0d737072
0000000a
65530a0d
5220646e
31313953
4c422e36
2e41542e
2e782e78
0d737072
0000000a
65530a0d
5220646e
31313953
4c422e36
2e344d2e
2e782e78
0d737072
0000000a
65530a0d
4b20646e
0a0d5945
00000000
65530a0d
4d20646e
0a0d5242
00000000
61530a0d
55206566
61726770
69206564
7250206e
6572676f
2e207373
0a0d2e2e
00000000
2059454b
61647055
53206574
65636375
75667373
000a0d6c
2052424d
61647055
53206574
65636375
75667373
000a0d6c
2059454b
61647055
46206574
656c6961
000a0d64
2052424d
61647055
46206574
656c6961
000a0d64
6f4c0a0d
6e696461
2e2e2e67
00000a0d
61560a0d
2064696c
6d726946
65726177
746f4e20
65725020
746e6573
00000a0d
6d490a0d
20656761
656e774f
694d2072
74616d73
0a0d6863
00000000
6c460a0d
20687361
20746f4e
65746544
64657463
00000a0d
6d490a0d
20656761
65746e49
74697267
61462079
64656c69
00000a0d
6f420a0d
4620746f
656c6961
000a0d64
70550a0d
64617267
6f697461
7553206e
73656363
6c756673
00000a0d
70550a0d
64617267
6f697461
7553206e
73656363
6c756673
44202620
75616665
4920746c
6567616d
766e4920
64696c61
7079422c
20737361
61736944
64656c62
00000000
70550a0d
64617267
6f697461
6146206e
64656c69
6552202c
7275422d
6874206e
6d492065
0d656761
0000000a
70550a0d
64617267
6f697461
6146206e
64656c69
646e6120
66654420
746c7561
616d4920
49206567
6c61766e
202c6469
61707942
44207373
62617369
0d64656c
0000000a
6e490a0d
696c6176
64412064
73657264
000a0d73
6f430a0d
6769666e
74617275
206e6f69
65766153
2e2e2e64
00000000
65440a0d
6c756166
6d492074
20656761
61766e49
0064696c
65440a0d
6c756166
6d492074
20656761
696c6156
00000064
52430a0d
61502043
64657373
00000000
52430a0d
61462043
64656c69
00000000
65440a0d
20677562
20676f4c
0000003a
0001c838
0001c854
0001bff0
00018004
0001ceef
0001cef0
614c0a0d
43207473
69666e6f
61727567
6e6f6974
746f4e20
76615320
00006465
6f420a0d
7075746f
74704f20
736e6f69
43524320
69614620
0064656c
45570a0d
4d4f434c
4f542045
44455220
454e4950
47495320
534c414e
00000000
6f420a0d
6f4c746f
72656461
72655620
6e6f6973
302e3120
0000302e
00000a0d
20310a0d
64616f4c
66654420
746c7561
72695720
73656c65
69462073
61776d72
00006572
20410a0d
64616f4c
72695720
73656c65
69462073
61776d72
28206572
67616d49
6f4e2065
30203a20
0029662d
20420a0d
6e727542
72695720
73656c65
69462073
61776d72
28206572
67616d49
6f4e2065
30203a20
0029662d
20350a0d
656c6553
44207463
75616665
5720746c
6c657269
20737365
6d726946
65726177
6d492820
20656761
3a206f4e
662d3020
00000029
204b0a0d
63656843
6957206b
656c6572
46207373
776d7269
20657261
65746e49
74697267
49282079
6567616d
206f4e20
2d30203a
00002966
20320a0d
64616f4c
66654420
746c7561
20344d20
6d726946
65726177
00000000
20330a0d
64616f4c
20344d20
6d726946
65726177
6d492820
20656761
3a206f4e
662d3120
00000029
20340a0d
6e727542
20344d20
6d726946
65726177
6d492820
20656761
3a206f4e
662d3120
00000029
20360a0d
656c6553
44207463
75616665
4d20746c
69462034
61776d72
28206572
67616d49
6f4e2065
31203a20
0029662d
20390a0d
63656843
344d206b
72694620
7261776d
6e492065
72676574
20797469
616d4928
4e206567
203a206f
29662d31
00000000
20460a0d
656c6553
4d207463
6e612034
69572064
656c6572
49207373
6567616d
61502073
00207269
20370a0d
62616e45
4720656c
204f4950
65736142
79422064
73736170
646f4d20
00000065
20380a0d
61736944
20656c62
4f495047
73614220
42206465
73617079
6f4d2073
00006564
20510a0d
61647055
4b206574
00005945
205a0a0d
4741544a
6c655320
69746365
00006e6f
20430a0d
6f636552
7269666e
6974616d
45206e6f
6c62616e
00000065
20440a0d
6f636552
7269666e
6974616d
44206e6f
62617369
0000656c
20480a0d
616e6942
4d207972
2065646f
62616e45
0000656c
20550a0d
616e6942
4d207972
2065646f
61736944
00656c62
20570a0d
73617245
69572065
656c6572
46207373
776d7269
20657261
616d4928
4e206567
203a206f
29662d30
00000000
20530a0d
73617245
344d2065
72694620
7261776d
49282065
6567616d
206f4e20
2d31203a
00002966
20260a0d
61647055
57206574
6c657269
20737365
0052424d
202a0a0d
61647055
4d206574
424d2034
00000052
6e450a0d
20726574
65726957
7373656c
616d4920
4e206567
2d30286f
0a0d2966
00000000
6e450a0d
20726574
4920344d
6567616d
286f4e20
29662d31
00000a0d
6e450a0d
20726574
4920344d
6567616d
69615020
6f4e2072
662d3128
200a0d29
0d20726f
0000000a
6e450a0d
20726574
6f742030
506e5520
0d726961
0000000a
6e450a0d
20726574
4741544a
74704f20
0d6e6f69
0000000a
6e450a0d
20726574
4f495047
6c655320
69746365
0a0d6e6f
00000000
65530a0d
7463656c
736f4820
300a0d74
52415520
310a0d54
49445320
320a0d4f
49505320
20340a0d
0d425355
5520350a
432d4253
0a0d4344
00000000
55200a0d
61726770
69746164
44206e6f
62617369
2c64656c
72754220
676e696e
20736920
20746f4e
6f6c6c41
2e646577
0a0d2e2e
00000000
6e450a0d
20726574
7478654e
6d6f4320
646e616d
00000a0d
61570a0d
7420746e
6843206f
65676e61
65687420
6e6f4320
75676966
69746172
203f6e6f
53455928
294f4e2f
000a0d20
6f430a0d
6769666e
74617275
206e6f69
6f6d6e55
69666964
2e2e6465
000a0d2e
61570a0d
6e697469
6f662067
6f432072
63657272
704f2074
6e6f6974
0d2e2e2e
0000000a
4d200a0d
6d492034
20656761
626d754e
49207265
6c61766e
0a0d6469
00000000
6e490a0d
696c6176
704f2064
6e6f6974
00000a0d
61560a0d
2064696c
6d726966
65726177
746f6e20
65727020
746e6573
00000a0d
00000004
0000000c
00000010
0000000c
00000014
00000018
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00101398
00101404
00101470
00101710
00101758
001018f4
00101824
00101880
00101990
00101a84
00101a34
00101dec
001050d0
00101e40
00101f00
001021b4
001022c8
001023cc
00103dac
001025f8
00102f00
00103450
001034c8
00103f4c
00103f70
0010401c
00104184
00104294
00104efc
00104924
00104860
001044b8
0010461c
00104318
001009b4
00100a00
001009d8
00102020
001051a4
001051d0
001051ec
0010522c
0010526c
00105294
001052bc
001052d4
00105308
00105388
001053c4
001053f4
0010541c
00105450
00105484
001054ec
00105554
00105724
001062b4
00105af0
00106034
00106068
00106368
001063a8
0010648c
001064b4
0010b900
0010b968
0010ba18
00100920
00100970
001011b0
001011dc
0010aaf4
0010ab3c
0010aee8
0010af4c
0010b5fc
0010b798
001009ac
00100f9c
00100d30
00100dc4
00100e8c
00100eb0
00100ee4
00100f70
00100f94
00106584
001065b8
001065dc
00106690
00114918
00114960
001149d8
00114a08
00114a34
0010bb58
00107ca0
0010bd7c
0010bc6c
00107974
00108944
0010bb9c
0010a340
0010a358
0010a368
0010a37c
0010a384
0010a38c
0010a394
0010a3a4
0010a3b4
0010a3c8
0010a414
0010a42c
0010a450
0010a530
0010a1fc
0010a234
0010a250
0010a25c
0010a280
0010a2a0
0010a2c8
0010a2f0
0010a318
0011103c
001066a0
001066c8
00106748
00106920
00106954
00106a1c
00106a84
00106aa4
00106aa8
00106b70
00106b80
00106c10
00106c40
00106c64
00106ca0
00106d10
00107a0c
00108004
00108030
001081fc
00108210
0010826c
001083a8
00108608
001088b8
0010a128
001091a4
00108f5c
00108ba0
00108ddc
0010960c
0010a01c
00100d00
00108cec
00108cb0
00108c78
0010958c
001089ec
0010897c
0010bc1c
001011fc
00101218
0010134c
001012f4
001122bc
001196c8
00119738
00119760
001197d4
00106558
0014d868
0014d8a0
0010aa70
0014d948
0014d9e8
0014dadc
0014db40
0014dd94
0014df40
001639e8
00157c5c
00163b78
00163b54
00163b34
00163ab8
00163a94
00163a74
00163b18
00163af4
00163ad4
00156b28
001638b4
00154a64
0015c630
0015e4c0
0015c9d0
0010a7b4
0010a808
0010a840
0010a958
0010a794
0010669c
00117868
001177d4
00117794
0011778c
001176a0
001178d8
00118394
001182e8
001181fc
0011850c
00118438
00117e5c
00117e50
001181bc
00118124
001180cc
00117e08
00118078
00118544
0011874c
00117944
00117998
001179a4
00117aa4
0010c6e8
0010c344
00118c68
00118cbc
0010c214
0011a8d0
001176d4
001173b0
001172ec
0011a374
0011a44c
0011a878
001175f4
001175d0
0011754c
00117408
00117414
0011742c
00117444
0011750c
00117454
001170c4
00116fc4
00116fcc
00118d64
001171c4
00100a44
00108e3c
001066dc
0010c2ec
00106e7c
0010b5bc
001075dc
00103484
0010a0d0
00112a84
00112b00
001085c0
0010bae4
0010d69c
0003e000
00437a31
40020000
00220000
007800d8
002000c7
00050001
00000000
00112ba0
00112bc4
00112c00
00112e1c
00112ea4
0011301c
0011306c
0011336c
001134d0
00113710
0011393c
00113b74
00113c00
00113d14
00114140
00114344
001144e4
00114918
00000000
00000000
0010a0d0
00113468
00114960
001149d8
00114a08
00114a34
001133c0
00114b5c
001140f0
00114c24
00114cb0
00114d20
001130e4
001130b0
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
00000000
40c31016
1341305c
201c6412
211c0dbc
0d000000
08729abc
345c7fe6
345c0ae7
345c0b27
08560b07
00000804
211c4046
680b4114
0100341c
2ef27df2
211c4306
680c4105
680f6092
211c4006
680b4114
5fff341c
63060253
4105311c
40724c0c
0dd24c0f
211c4006
680b4114
7fff341c
680b680e
6d723364
0153680e
311c6006
4c0b4114
a000101c
236421a3
08044c0e
0136f016
71c340c3
53c362c3
0b84801c
0000811c
0004f524
00040004
706c502c
702f32a3
506f4006
c5f20433
0004f324
00040004
08ce0cbc
0a1d373c
001c67d2
011c0bb4
36640000
011600f3
680c28c3
36640e86
c0278056
f3240594
00040004
f5240004
00040004
500c0004
704c102c
03830283
da940007
102c300c
704c506c
20a33183
66d23283
0004f324
00040004
a3f2f853
f7f31404
f7b35664
0f568076
00000804
200f2006
402f5fe6
206f404f
00000804
8e243016
213cf524
301c200c
311c0fe4
ac0c0000
440c2a80
30236026
640f32a3
4004343c
f32462d2
08040c56
8e241016
213cf524
301c200c
311c0fe4
2c0c0000
280c4880
30236026
318333e3
343c680f
62d24004
0856f324
00000804
8e241016
213cf524
301c200c
311c0fe4
2c0c0000
282c4880
30236026
318333e3
343c682f
62d24004
0856f324
00000804
8e241016
213cf524
301c200c
311c0fe4
2c0c0000
284c4880
30236026
318333e3
343c684f
62d24004
0856f324
00000804
8e243016
213cf524
301c200c
311c0fe4
ac0c0000
442c2a80
30236026
642f32a3
4004343c
f32462d2
08040c56
8e243016
213cf524
301c200c
311c0fe4
ac0c0000
444c2a80
30236026
644f32a3
4004343c
f32462d2
08040c56
40c33016
f524ae24
200c213c
0fe4301c
0000311c
28000c0c
6026042c
400d233c
308332e3
646c642f
446f23a3
4004353c
f32462d2
08040c56
200c213c
0fe4301c
0000311c
68802c0c
033c6c0c
041c008d
08040001
200c213c
0fe4301c
0000311c
68802c0c
6c4c4c0c
30833283
602662d2
080403c3
200c213c
0fe4301c
0000311c
68802c0c
033c6c2c
041c008d
08040001
31c31016
f5242e24
200c233c
0fe4301c
0000311c
6a008c0c
313c0c4f
62d24004
0856f324
00000804
31c31016
f5242e24
200c233c
0fe4301c
0000311c
4a008c0c
03a3684c
313c084f
62d24004
0856f324
00000804
8e243016
213cf524
301c200c
311c0fe4
ac0c0000
444c2a80
328330e3
343c644f
62d24004
0c56f324
00000804
50c37016
ce2441c3
648bf524
0b1403e4
301c0116
311c0b84
6c0c0000
009f001c
80563664
35236026
502c33e3
702f3283
10ab64f2
089570bc
4004363c
f32462d2
08040e56
40c37016
ce2451c3
8ebcf524
740c0895
4e1d333c
00070c20
60260674
542c3423
62f23283
363c0006
62d24004
0e56f324
00000804
1f36f016
61c390c3
b1c32e24
982cf524
0001a01c
8ebc04d3
80c30895
0cbc04c3
10c308ce
000d3a3c
182c73e3
60073083
513c1754
580c180c
1e1d323c
feb0c33c
301cc8a4
311cffea
83c37fff
0835c8e4
308337c3
6a80782f
09c36c2c
47833664
da948007
08958ebc
982c70c3
801cbfe6
02730001
0cbc04c3
780c08ce
0e1d333c
40074fa0
a0860315
383c0153
33e3000d
52e44383
52c30235
ed948007
6007782c
a2f21354
38aba026
341c31c3
201c000f
211c0fe4
494c0000
200603c3
5000111c
15c301a3
3b3c2664
62d24004
f876f324
08040f56
0736f016
91c360c3
2e2453c3
f524a1c3
600672c3
8000311c
42c37383
748b9f92
0b1443e4
301c0116
311c0b84
6c0c0000
009f001c
80563664
c007edf2
01160b15
0b84301c
0000311c
001c6c0c
3664009e
60268056
400d833c
342c38e3
742f3183
08958ebc
06c310c3
0700e2f2
180c343c
6d00540c
740c2c31
4f9d033c
800780a0
802602d4
14ab742c
303c64f2
019300f4
089580bc
143440e4
62676220
54ab1135
341c32c3
201c000f
211c0fe4
494c0000
200603c3
5000111c
14c301a3
742c2664
742f38a3
40043a3c
f32462d2
0f56e076
00000804
0136f016
71c340c3
63c352c3
82c34e24
05c3f524
13c31f92
0873d6bc
073404e4
17c304c3
36c325c3
08745abc
4004383c
f32462d2
0f568076
00000804
60c37016
200702c3
51c31d54
53837f86
800602c3
7a0100f3
03e40180
00250234
45e48085
141cf914
2cd20003
180c213c
32237fe6
5a0133e3
0c003283
023403e4
0e560025
00000804
70c3f016
52c361c3
42c34006
073c0133
163c4a1d
e2bc4a1d
20c30874
45e48025
02e3f714
08040f56
311c6006
201c4113
4c0e0150
311c6006
201c4008
4c0e1150
00000804
4ccc604c
0204301c
4130311c
32c34c0f
305c6492
08040427
60c37016
0218301c
4130311c
00062c0c
00ff011c
401c1083
411c0210
b00c4130
00064c0c
00ff011c
21e42083
12c30334
301cfef3
311c0084
6c0b4040
436443c3
011c0a06
600c4140
000f341c
64d22026
133c600c
503200f4
3410141d
3230141d
780f6e80
08040e56
60c3f016
0218301c
4130311c
00062c0c
00ff011c
401c1083
411c0210
b00c4130
4c0cf02c
011c0006
208300ff
033421e4
fed312c3
0084301c
4040311c
43c36c0b
0a064364
4140011c
341c600c
2026000f
600c64d2
00f4133c
141d5032
141d3410
6e803230
4006780f
023435e4
6b804026
0f56782f
00000804
41c33016
13c352c3
341c30c3
6dd23fff
708c203c
32236026
32a3440c
021c640f
301c4000
0383c000
341c34c3
6bd23fff
708c243c
32236026
32a3440c
301c640f
4383c000
113404e4
133c7020
4026708c
303c0173
323c708c
940c300d
740f34a3
4000021c
36f23fe5
08040c56
211c42c6
680b4105
66723364
301c680e
311c0880
40062200
60854c0f
0100201c
61054c0f
00f8201c
301c4c0f
311c0888
201c2200
4c0f03c6
0361305c
61cc64f2
36646e0c
00000804
0200301c
4130311c
4c0f4026
00000804
211c49c6
680b2100
0004341c
608666d2
6006680e
05a7305c
00000804
83c61016
2100411c
341c700b
67d20004
6d4c616c
60863664
0073700e
10041004
08040856
0736f016
71c340c3
93c382c3
af5ca257
603c0144
305c1640
602705a4
01160b94
0b84301c
0000311c
001c6c0c
366400b2
00068056
031550e4
0086bf92
245c4006
745c0b87
63970b27
fc2c333c
0b47345c
0016353c
0b0d333c
233c7fe5
6217f88c
d1ac393c
3a3c6e72
3a3ca1ac
323c81ac
345c79ac
26c30b67
301c2364
311c0098
4c0e2100
808c263c
4c0e6045
f5242e24
0b0d353c
233c7fe5
303cf88c
223c0815
694659ac
2100311c
60264c0e
05a7345c
4004313c
f32462d2
0f56e076
00000804
05a4305c
30546007
211c49c6
20072100
4e241e54
29c6f524
2100111c
341c640b
64f20004
05a4305c
69c66af2
2100311c
2c0e2086
4004323c
02d368f2
f5241404
00040004
fd730004
01d3f324
341c680b
65f20004
341c680b
79f20001
311c69c6
40862100
60064c0e
05a7305c
00000804
0736f016
51c340c3
83c362c3
0104af5c
01249f5c
1640703c
05a4305c
0b946027
301c0116
311c0b84
6c0c0000
00b2001c
80563664
345c6006
545c0b87
645c0b27
3a3c0b47
333c0016
7fe50b0d
f88c233c
6e7238c3
a1ac393c
81ac393c
79ac323c
0b67345c
236427c3
0098301c
2100311c
273c4c0e
6045808c
2e244c0e
201cf524
3ac30881
201c63d2
69460081
2100311c
40264c0e
05a7245c
4004313c
f32462d2
0f56e076
00000804
05a4305c
11546007
211c49c6
680b2100
0004341c
680b65f2
0001341c
69c679f2
2100311c
4c0e4086
305c6006
080405a7
ff96f016
203740c3
7f5c63c3
5f5c00c3
31c30001
0400341c
ffff001c
020f011c
60073400
313c1054
133c200c
640b00e0
0004341c
640b65f2
0001341c
608679f2
0173640e
200c313c
6c0b61c5
0001341c
60070026
000854dc
106f0006
d02f500f
304f21d7
32c34017
0100341c
fff0053c
101c6bd2
111c00dc
440b2100
30236026
336432a3
101c0173
111c00dc
440b2100
60262364
33e33023
640e3283
30c30017
0200341c
0070053c
101c6bd2
111c00dc
440b2100
30236026
336432a3
101c0173
111c00dc
440b2100
60262364
33e33023
640e3283
0067153c
311c6f46
45802100
336434c3
0f86680e
2100011c
343c4400
680e808c
ffff101c
020f111c
133c7480
213c200c
37c300a0
680e6272
32c34017
0800341c
23546007
341c32c3
213c1000
600700e0
4e241654
21c5f524
341c640b
67d20004
640e6086
4004323c
01f368f2
f5241404
00040004
fe330004
00f3f324
341c680b
7dd20004
080e0086
01960006
08040f56
40c33016
211c41c6
680b2100
0004341c
31546007
680e6086
6007632c
301c2894
311c0bb4
535c0000
744c0764
11946007
01dc021c
c710101c
0011111c
44bc4086
01640892
0b0d303c
7f3233c4
744f6025
0ee4145c
28d2716c
04c36ccc
60063664
0ee7345c
6d0c0153
007304c3
6d0c616c
00733664
10041004
08040c56
0336f016
90c3fe96
61c373c3
341c31c4
49a00003
3c0900b3
c02561c3
7cf27fe5
0034023c
30c33900
9c090093
7fe5840d
7cf23fe5
6257a820
d005833c
45c30373
1f00531c
401c0335
201c1f00
40370081
341c34c3
101c1fff
111c4000
31a30110
09c36077
27c318c3
2abc36c3
b6200877
a007da00
0296e594
0f56c076
00000804
211c4006
680c4140
680f7072
680c4705
680f7972
00000804
211c4006
680c4140
680f7092
680c4705
680f7992
00000804
fd963016
126453c3
20278306
83860554
02542047
64068406
412c311c
1000001c
60450c0e
133c6c0b
1fe61004
3b942007
311c6486
02a6412c
00060c0e
412c011c
6c0b6400
013c68c1
00b70020
00411f5c
f41414e4
311c6486
02c6412c
40060c0e
111c2006
6880412c
75416c0b
0020023c
2f5c0077
24e40021
6486f414
412c311c
4c0e42e6
00064006
412c011c
6c0b6800
65412197
0020023c
2f5c0037
24e40001
0006f314
0c560396
00000804
fb96f016
72c361c3
026453c3
44060137
412c211c
0080001c
8306080e
21176006
002701c3
83860c54
0400301c
01c32117
05540047
280e2806
60068406
036403c3
0055303c
236423c3
311c6486
4c0e412c
40062006
412c211c
58e26500
213c4c0e
40f70020
00611f5c
f41414e4
0065303c
236423c3
311c6486
4c0e412c
40062006
412c211c
5ce26500
213c4c0e
40b70020
00411f5c
f41414e4
0075303c
236423c3
311c6486
4c0e412c
00062006
412c011c
54e26400
313c4c0e
60770020
00211f5c
f41414e4
311c6406
4c0b412c
43722364
44464c0e
412c211c
341c680b
7dd20008
0066a037
00812f5c
26c312c3
72bc37c3
05960878
08040f56
3f36f016
83c3f996
0304bf5c
0324cf5c
0344df5c
01b70264
526451c3
626462c3
02a17f5c
02c1af5c
02e19f5c
08785abc
311c6406
001c412c
0c0e0080
20068306
02c34197
12540027
101c8386
41970400
004702c3
80060b54
419714c3
008702c3
28060594
84062c0e
a0072006
44c66f54
412c211c
680e6026
680bc5d2
62723364
0197680e
64c608f2
412c311c
23644c0b
00f34372
311c64c6
4c0b412c
44722364
a0474c0e
64863294
412c311c
ac0ea1c6
211c4006
0197412c
14940007
c718501c
0011511c
00066a80
bed4011c
6c0b6c00
016f323c
311c6a46
53c3412c
ef9425e4
001c06b3
011cc730
68000011
511ca006
6e80bed4
323c6c0b
0ec6016f
412c011c
23e430c3
0453ef94
2094a027
311c6486
41c6412c
60064c0e
412c311c
6045ac0e
abf2a197
033c0006
4a46016f
412c211c
35e452c3
0153f894
033c0006
4ec6016f
412c211c
35e452c3
01c3f894
64860364
412c311c
20060c0e
400601b3
412c211c
58c36500
4c0e54e2
0020313c
1f5c6177
14e400a1
30c3f314
23c36172
64862364
412c311c
20064c0e
400601b3
412c211c
a4976500
4c0e54e2
0020313c
1f5c6137
14e40081
303cf314
23c30035
64862364
412c311c
20064c0e
400601b3
412c211c
a4d76500
4c0e54e2
0020313c
1f5c60f7
14e40061
30c3f314
23c36272
64862364
412c311c
17c34c0e
2254e007
311c6006
0026412c
40460c0e
20060193
412c111c
a0066880
123cac0e
20b70020
00412f5c
f41424e4
a0060813
412c511c
05176680
4c0e40e2
0020313c
1f5c6077
14e40021
09c3f314
640608d2
412c311c
23644c0b
4c0e4872
311c6406
4c0b412c
40722364
19c34c0e
27942007
211c4446
680b412c
0001341c
df5c7dd2
00060007
00c12f5c
2bc312c3
72bc3cc3
3ac30878
5f5c69d2
05c300c1
2cc31bc3
c8bc3dc3
66bc0878
01330878
311c6406
4c0b412c
44722364
f9134c0e
fc760796
08040f56
3f36f016
62c3f696
bf5c73c3
cf5c0384
df5c03a4
026403c4
91c30277
5f5c9264
af5c0321
8f5c0341
5abc0361
44060878
412c211c
0080301c
0306680e
82576006
202714c3
03860c54
0400301c
14c38257
05542047
680e6806
60060406
436443c3
0055343c
236423c3
311c6486
4c0e412c
40062006
412c211c
58e26500
213c4c0e
42370020
01011f5c
f41410e4
0065343c
236423c3
311c6486
4c0e412c
c0062006
412c611c
5ce26700
313c4c0e
61f70020
00e11f5c
f41410e4
0075343c
236423c3
311c6486
4c0e412c
a00715c3
60061554
412c311c
2c0e2026
c0064046
412c611c
20066b00
623c2c0e
c1b70020
00c12f5c
f41420e4
400601f3
412c211c
c5576500
4c0e58e2
0020313c
1f5c6177
10e400a1
34c3f314
23c36172
64862364
412c311c
20064c0e
211c4006
6500412c
58e2c597
313c4c0e
61370020
00811f5c
f31410e4
0035343c
236423c3
311c6486
4c0e412c
40062006
412c211c
c5d76500
4c0e58e2
0020313c
1f5c60f7
10e40061
34c3f314
23c36272
64862364
412c311c
15c34c0e
1554a007
311c6006
2026412c
40462c0e
411c8006
6a00412c
cc0ec006
0020323c
2f5c60b7
20e40041
0933f414
611cc006
6700412c
50e28617
213c4c0e
40770020
00211f5c
f31410e4
88d248c3
311c6406
4c0b412c
4a722364
69c34c0e
6486c8d2
412c311c
23644c0b
4c0e4872
311c6406
4c0b412c
42722364
18c34c0e
27942007
211c4446
680b412c
0004341c
df5c7dd2
00260007
01212f5c
2bc312c3
72bc3cc3
3ac30878
4f5c69d2
04c30121
2cc31bc3
c8bc3dc3
66bc0878
01330878
311c6406
4c0b412c
44722364
f7f34c0e
fc760a96
08040f56
0136f016
51c3fb96
83c372c3
01370264
01616f5c
08785abc
211c4406
001c412c
080e0080
60068306
01c32117
0c540027
301c8386
21170400
004701c3
28060554
8406280e
03c36006
303c0364
23c30055
64862364
412c311c
20064c0e
211c4006
6500412c
4c0e54e2
0020213c
1f5c40f7
14e40061
303cf414
23c30065
64862364
412c311c
20064c0e
211c4006
6500412c
4c0e5ce2
0020213c
1f5c40b7
14e40041
303cf414
23c30075
64862364
412c311c
20064c0e
011c0006
6400412c
40e208c3
313c4c0e
60770020
00211f5c
f31414e4
6406c8d2
412c311c
23644c0b
4c0e4972
311c6406
4c0b412c
41722364
c0074c0e
44461494
412c211c
341c680b
7dd20002
20372397
2f5c0046
12c30081
63574317
087872bc
087866bc
80760596
08040f56
ff967016
126450c3
211c4486
60062040
313c680e
351c480c
33640009
0206680e
030625d2
02542027
40060406
411c8506
28062040
2040111c
341c700b
7df20004
640f7501
0040623c
2f5cc037
20e40001
4506f414
2040211c
341c680b
7dd20001
0e560196
00000804
313c1016
341c480c
233cfe00
64860115
2040311c
40064c0e
411c8506
28062040
2040111c
341c700b
7df20004
640f6101
42074085
4506f894
2040211c
341c680b
7dd20001
08040856
6586200c
2040311c
202c2c0f
2c0f6085
6085204c
406c2c0f
4c0f6085
00000804
0136f016
70c3f896
226481c3
126413c3
01c13f5c
43f26912
00736072
0005351c
236423c3
311c6486
4c0e2040
08942027
311c6486
4c0b2040
41722364
20470133
64860894
2040311c
23644c0b
4c0e4672
10fc601c
0000611c
6cc9780c
2b946007
850613c3
2040411c
611cc806
a8862040
2040511c
400603b3
700b1c80
0004341c
61017df2
4085780f
f8944207
341c700b
7dd20001
63d74006
700b0c80
0020341c
740c7df2
40856161
f8944207
18e42205
0cf3e314
01004f3c
220604c3
08cb9cbc
22060fc3
08cb9cbc
311c6406
22262040
e1372c0e
211c4806
4177a040
001c38c3
011c4000
30a30001
288661b7
a040111c
43d72037
60b74077
cd29780c
103c0d09
6f460067
2100311c
34c34580
680e3364
311c6f86
45802100
808c343c
163c680e
6f460067
2100311c
3fc34580
680e3364
311c6f86
45802100
808c3f3c
101c680e
111cffff
6080020f
200c233c
00a0323c
0085001c
78800c0e
200c133c
00a0313c
41c50c0e
341c680b
7dd20004
680e6086
00e0213c
341c680b
7dd20004
080e0086
311c6486
20062040
08962c0e
0f568076
00000804
0f36f016
a0c3f996
72c351c3
83c37264
4f5c8264
4e240201
f524b2c3
78bc0126
673c08cc
c0b7ffd0
00411f5c
926491c3
0080601c
0001931c
c8060235
600738c3
301c7294
311c0200
4c0c2040
4c0f4772
0204201c
2040211c
341c680c
7dd20200
0200301c
2040311c
273c4c0c
4c0f192c
10b4e047
6105540c
542c4c0f
4c0f6105
6105544c
546c4c0f
4c0f6105
6105548c
373c4c0f
6077fff0
00213f5c
0db46027
301c54ac
311c0230
4c0f2040
610554cc
54ec4c0f
4c0f6105
0001931c
540c3cb4
0208301c
2040311c
542c4c0f
4c0f6085
6085544c
546c4c0f
4c0f6085
6085548c
54ac4c0f
4c0f6085
608554cc
54ec4c0f
4c0f6085
6085550c
552c4c0f
4c0f6085
6085554c
556c4c0f
4c0f6085
6085558c
55ac4c0f
4c0f6085
608555cc
55ec4c0f
01136085
0200301c
2040311c
273c4c0c
4c0f192c
0200301c
2040311c
42724c0c
80074c0f
163c1894
24c3108c
0204401c
2040411c
0280001c
2040011c
341c700c
7df20080
363c6ac3
600f2a1d
21e44025
07b3f614
00c04f3c
220604c3
08cb9cbc
0067af5c
0280101c
2040111c
201c2137
211c4000
62a30c01
301cc177
311c10fc
6c0c0000
103c0ce9
6f460067
2100311c
34c34580
680e3364
611ccf86
47002100
808c343c
101c680e
111cffff
6080020f
200c233c
00a0323c
0085601c
41c5cc0e
341c680b
7dd20004
280e2086
fff0383c
f88c033c
831c05f2
44dc0002
101c000b
111c0204
640c2040
1004233c
301c5df2
311c0200
4c0f2040
0204201c
2040211c
341c680c
7dd20001
0208301c
2040311c
740f6c0c
0001931c
301c5bb4
311c020c
6c0c2040
301c742f
311c0210
6c0c2040
301c744f
311c0214
6c0c2040
301c746f
311c0218
6c0c2040
301c748f
311c021c
6c0c2040
301c74af
311c0220
6c0c2040
301c74cf
311c0224
6c0c2040
301c74ef
311c0228
6c0c2040
301c750f
311c022c
6c0c2040
301c752f
311c0230
6c0c2040
301c754f
311c0234
6c0c2040
301c756f
311c0238
6c0c2040
301c758f
311c023c
6c0c2040
301c75af
311c0240
6c0c2040
301c75cf
311c0244
6c0c2040
e04775ef
301c19b4
311c0210
6c0c2040
301c742f
311c0218
6c0c2040
301c744f
311c0220
6c0c2040
301c746f
311c0228
6c0c2040
273c748f
4037fff0
00013f5c
13b46027
0230301c
2040311c
74af6c0c
0238301c
2040311c
74cf6c0c
0240301c
2040311c
74ef6c0c
301c07d2
311c0200
20062040
01262c0f
08cc82bc
40043b3c
f32462d2
07960006
0f56f076
00000804
0bb4301c
0000311c
2c4c4cec
03c348ac
26642b05
00000804
0bb4301c
0000311c
2c4c4cec
03c348ac
0098121c
08042664
6027646c
642c1594
12946087
0c44305c
301c68d2
311c0100
4c0c4130
00f34f72
00a4301c
4140311c
43724c0c
08044c0f
65ac000c
0074133c
606c25f2
06e4335c
08043664
60c3f016
e04c51c3
341c7c8c
60070002
620c2854
36646e0c
341c75ac
60070007
301c1194
311c801c
101c4113
2c0e5400
4000301c
4128311c
803b201c
0000211c
301c01d3
311c801c
101c4113
2c0e5000
4000301c
4128311c
01a0201c
02f34c0f
55ec206c
190b323c
153c840c
241c03d0
4664000f
341c75ec
69d20008
8c2c786c
04c0053c
255c13c3
46640303
211c4006
680b4008
dfff341c
766c680e
0020341c
1b546007
6c4c78ec
15c306c3
55ac3664
0784323c
08546f07
6d8c78cc
15c306c3
09cb223c
7c8c3664
0002341c
78ec66d2
06c36c8c
366415c3
61927c8c
0f567c8f
00000804
40c37016
c0eca04c
63f276ac
64d2762c
04c3792c
766c3664
722c65d2
04c36c6c
