09f8eebc
104d0264
306d2006
4546f02f
312d510d
00d4055c
f8bc19c3
b64b09f7
3f5ca137
714d0081
08320117
1f5c00f7
316d0061
40c60433
6006500d
06c3702d
09f8eebc
104d0264
106d0006
27c6f02f
112d310d
153c09c3
42060160
08cbb0bc
a077b78b
00212f5c
6057514d
60376832
00010f5c
1ac3116d
6a0c440c
6a0f6025
01592f5c
323c4277
1bc303c7
4f496580
341c32c3
60070008
301c1054
311c1110
6c0c0000
0544335c
01211f5c
18c301c3
30c33664
6bf23264
1110301c
0000311c
335c6c0c
00060484
366418c3
f0760d96
08040f56
0736f016
81c370c3
536452c3
202ba0c3
28c3a184
301c4af2
311c0b84
6c0c0000
2454001c
07933664
a3f2c006
01f365c3
180c363c
2ccb7d80
091451e4
53c374a0
363c5364
63c30010
b3f26364
0293975c
cef204b3
44891ac3
620532c3
08c36e80
7ccb2580
b0bc4ea0
3ccb08cb
263c0213
363c0010
9d80180c
373c08c3
35802e1d
063e343c
b0bc4ea0
300b08cb
838466a0
0010363c
636463c3
69e4a006
e076db14
08040f56
fe961016
616c40c3
202640cc
00061f5c
1f5c2006
00060025
30c313c3
0a79b2bc
408c0cd2
313c318b
638e0100
313c680c
680f601b
684d6026
08560296
00000804
ff967016
301c60c3
311c1110
6c0c0000
0af28c0c
0b84301c
0000311c
001c6c0c
36642456
503c0b13
748cf680
2037200c
07942027
00011f5c
40462c4d
05934c8d
13c36017
14942047
0a00bcbc
000750c3
500c2394
6025688c
301c688f
311c0bb4
0c0c0000
25c316c3
08e6e6bc
bcbc0693
50c30a00
796c0bf2
796f61c5
7e4578cc
06c378cf
0a0ae8bc
780c04d3
700c65f2
40254ccc
784c4ccf
aaaa201c
aaaa211c
31e412c3
7fe70654
60260454
04a7355c
0cbc05c3
8e240a05
301cf524
311c1110
6c0c0000
06c36f2c
366415c3
4004343c
f32462d2
0e560196
00000804
3f36f016
60c3fa96
326431c3
00066077
301c0177
311c1110
6c0c0000
301cec0c
311c0bb4
4c100000
01c1175c
7c0c26f2
40254dcc
31b34dcf
582b96c3
a0069284
535c39c3
b35c002e
3b3c0021
89c30100
d65c8384
c65c0003
18c30013
32c345a9
12c34589
41ac413c
533c38c3
03c3071e
09f812bc
00f70364
8066343c
fff0233c
361c34c3
7fe58035
033c32a3
00b7f88c
21372086
353c04f2
6137208c
35c3a117
0006361c
133c7fe5
2037f88c
40d726d2
658732c3
0014e2dc
a9d2a017
05067dec
0002011c
60073083
001442dc
ff003d3c
3ba43ca4
b364b3c3
14c308c3
23c360d7
00815f5c
70bc35c3
10c309f8
5c0c1264
42dc2007
698c0013
698f6025
10c30117
a4dc2087
07330009
6e2c6c0c
009340c6
6e2c6c0c
36644086
59c34157
182bb489
62057400
692f7980
582b2157
59c332c4
6ea0b489
1f00233c
6d00652c
0097654f
431c0cf2
09540800
86dd201c
0000211c
43e432c3
000fe4dc
ad2c6157
6157ad6f
61576cd1
0ccc4d6c
4d8f4800
21571c4c
eabc4057
20b30a40
2fd22097
1f3c1d4c
44860140
5abc6006
00070a4e
000e24dc
4d6c6157
0fb35e45
0800431c
000974dc
53c360d7
2094a0c7
015c18c3
303c0174
6cf28004
210b303c
64456212
0454b3e4
003cb31c
1d4c03b4
1c6c0053
01401f3c
60064706
0a4e5abc
b4dc0007
6157000b
59454d6c
5f5c0ad3
35c30041
10c300d7
04942027
00612f5c
326432c3
05c3a0d7
06540227
25c365f2
08544047
66d21453
1f3c1d4c
48060140
1c6c00b3
01401f3c
60064586
0a4e5abc
34dc0007
61570009
5ac54d6c
601705d3
b2dc6007
501c0008
511c86dd
05c30000
389440e4
21c320d7
219440c7
035c38c3
403c0214
8df28004
210b303c
66c56212
0794b3e4
1f3c1d4c
49860140
00d334c3
1f3c1c6c
49860140
5abc6006
00070a4e
61576494
56c54d6c
03934d6f
01401f3c
20c300d7
03944747
00531d4c
48061c6c
5abc6006
61570a4e
58454d6c
0ad24d6f
301c0993
311c0b84
6c0c0000
2455001c
60d73664
a02753c3
b31c0494
08b4015e
21c320d7
0d944747
0172b31c
7c0c0a35
40254dec
01574def
0a4066bc
a177a006
40074157
694c2654
092c7fc5
b3e46c20
301c1915
311c1110
6c0c0000
04e4335c
296c06c3
36644006
6cd16157
4d6c6157
4a80accc
1c4c4d8f
40572157
0a40eabc
7c0c0113
40254dec
01574def
0a4066bc
4dac7c0c
4daf4025
16c30ac3
08e71abc
696c0293
696f6025
0580063c
301c0177
311c1110
201c0000
211c86dd
52c30000
b4dc45e4
d8b3ffec
fc760696
08040f56
fe961016
301c0364
311c1110
6c0c0000
303c4c0c
082c03c7
4c0c6c00
40074077
6e691f54
20772026
1a9460c7
025c2006
40c30201
0209025c
422c303c
0211425c
81ac343c
0219025c
c1ac303c
025460a7
413c2026
80370016
00010f5c
1f5c0077
01c30021
08560296
00000804
f8963016
600650c3
61b761f7
106c301c
0000311c
301c2c0c
311c1110
6c0c0000
4c4c6c0c
01803f3c
85ac6037
202602c3
00402f3c
01c03f3c
05c34664
00801f3c
b0bc4206
089608cb
08040c56
fe961016
126440c3
00770006
301c0037
311c1110
6c0c0000
6b0b4c0c
169460a7
0a942027
0229325c
04946027
01a1125c
000601d3
2af20273
0229325c
06946027
01a1025c
13c304f2
20060053
2f3c084c
3fc30040
0a625ebc
14c30057
09f7f8bc
08560296
00000804
1f36f016
70c3f096
1110301c
0000311c
2c106c0c
433c608c
30490100
a45c20f7
313c0019
19c303c7
cc80242c
41375a69
305c6006
20d704a7
0ebc01c3
30c30a03
60073264
784c4554
4c8964d2
40544007
13c37149
b33c7169
300940ac
302921c3
412c513c
1594a087
03800f3c
6abc3a49
3f5c0a03
600701c1
1f5c1b94
200701c9
2f5c1794
400701d1
3f5c1394
01d301d9
0e94a0c7
02800f3c
0a0344bc
68f26297
66f262d7
64f26317
60076357
41171154
60c732c3
786c1b94
18546007
a0876906
6b860254
69a05f8b
056e331c
301c0ff4
311c0ef0
4c0c0000
0bb4301c
0000311c
173c0c0c
26640040
143c1af3
a08700c0
a1771794
03c00f3c
b0bc25c3
3f5c08cb
701201e9
01e14f5c
c1ac343c
01f91f5c
2f5c31a3
323c01f1
61b741ac
60c60113
0f3c6177
42060180
08cbb0bc
6007784c
8c892d54
2a548007
1000073c
a087600c
341c0794
533c0fff
2706fc80
341c00d3
533c0fff
2986fb40
0006801c
0083531c
801c0335
301c0008
311c1110
4c0c0000
0100313c
60376180
0a3c89f0
2026388c
00f42a3c
762048c3
401cc664
411c1110
700c0000
07c36e0c
00812f5c
415712c3
50c33664
13c36117
1e942227
8e4c700c
15c3180c
01402f3c
46643bc3
0f5c0077
00070021
39c37354
682c4c0c
682f6025
700c49c3
301c0c0f
311c0b84
6c0c0000
448d001c
21170b13
40c721c3
ee245794
3a09f524
341c31c3
6bf20001
40075a4b
700c1a94
180c6eac
366415c3
13540007
1110301c
0000311c
6ecc6c0c
15c3180c
36644006
0f5c00b7
373c0041
60074004
02731394
4004373c
f32462d2
1110301c
0000311c
6fac6c0c
00614f5c
15c304c3
366429c3
f3240573
28540007
640c19c3
303c0c0f
7fe50396
63f27f32
0c940927
500c49c3
684c65d2
684f6025
686c01b3
686f6025
301c0133
311c0b84
6c0c0000
448e001c
1fe63664
301c0153
311c0b84
6c0c0000
248f001c
00063664
f8761096
08040f56
1110301c
0000311c
6c0c6c0c
033c6cec
080401d0
1110301c
0000311c
6c0c6c0c
033c6d0c
08040140
40c31016
1110301c
0000311c
680c4c0c
20066dec
1000111c
65d23183
00066b4c
366414c3
1110301c
0000311c
6f6c6c0c
366404c3
08040856
f5244e24
2344305c
323c69f2
62d24004
01c3f324
0a4066bc
305c03d3
241c22c4
6cd20400
22e4305c
60062c2f
105c642f
400722e7
f3241054
105c01d3
105c22c7
642f22e7
f32442d2
01fc021c
40062206
09e0bebc
00000804
40c3f016
63c352c3
36544007
001c680c
011c434b
20c35041
2e9432e4
2c548007
2a542007
0046716c
27c3f12c
271432e4
0066718c
27c3f14c
21b432e4
1654c007
11b4301c
0000311c
40074c0c
301c1754
311c139c
6c0c0000
10946007
12c0301c
0000311c
27e473c3
04c30954
36c325c3
0a0a06bc
00e60093
02260053
08040f56
0136f016
40c3ff96
53c362c3
6007e1d7
6c0c3a54
434b001c
5041011c
32e420c3
80073294
20073054
01262e54
2e54c007
0046716c
82c3512c
281438e4
0066718c
82c3514c
22b438e4
1654e007
11b4301c
0000311c
40074c0c
301c1854
311c139c
6c0c0000
11946007
12c0001c
0000011c
23e430c3
e0370a54
26c304c3
6ebc35c3
00930a0a
005300e6
01960226
0f568076
00000804
40c31016
600c000c
15356047
18546007
201c6c0c
211c434b
12c35041
109431e4
412c616c
31e412c3
618c0b14
12c3414c
06b431e4
0a4066bc
100f04f2
00e60053
08040856
40c31016
0007000c
600c1b54
18546007
101c6c0c
111c434b
21c35041
109432e4
212c616c
32e421c3
618c0b14
21c3214c
06b432e4
0a0ae8bc
100f04f2
00e60053
08040856
0736f016
70c3ff96
42c351c3
901c4710
801c0028
811c106c
d7ab0000
22dc8647
8647000e
856707b4
85874054
8bd25254
86670c73
000d72dc
42dc8767
8787000d
01b35b94
106c201c
0000211c
01c1355c
47946007
155c2026
047301c5
01c9355c
01c1255c
04946027
08b44027
40470173
204605b4
01c5155c
40e60093
01c5255c
155c6006
21c301c9
40374025
00011f5c
01cd155c
106c201c
0000211c
21946007
680c28c3
01f36dcc
01c1355c
106c201c
0000211c
15b46047
255c4066
18c301c5
6dec640c
15c307c3
00073664
11736a54
01c1355c
106c201c
0000211c
03356067
0ad3680c
355c6086
680c01c5
07c36e0c
366415c3
55ec0f13
0c9480c7
07544087
709440c7
68492ac3
6c946087
1b84375c
40c704b3
87470694
375c0494
03d315e4
0046323c
0b0d333c
7f327fe5
802766d2
375c0494
02531584
804766d2
375c0494
019314a4
11948227
40c767f2
1ac34b94
60876449
375c4794
60071904
07c34354
366415c3
07f30006
0964375c
07c369d2
800c143c
366425c3
600730c3
75ec3454
309460c7
106c301c
0000311c
8e2c6c0c
15c307c3
211c4006
36c30401
04534664
60c775ec
fff3b4dc
8409356c
86676429
62120594
0020233c
60250093
180c233c
62e4d4cc
00260334
650000b3
7920756f
955c74cf
556c01d6
04f2772c
93a492c3
0026e3b3
e0760196
08040f56
6e241016
205cf524
433c0924
4cd24004
0944305c
60062c2f
105c642f
80070947
f3241054
105c01d3
105c0927
442f0947
f32482d2
01fc021c
40062106
09e0bebc
08040856
64f264ec
4a80303c
456c64ef
64526808
472f65ef
04946087
2984305c
60c700b3
305c0694
63d23144
00933664
66bc01c3
08040a40
43c3f016
a00631c3
f000511c
c0063583
e000611c
37e476c3
3fe70354
300f0b94
6006280c
32942007
4a80303c
31c3680f
505c05b3
acd22561
4a80503c
605c31c3
36832604
2624705c
36e467c3
705c1054
e0072781
503c1154
31c34ec0
2824605c
705c3683
67c32844
069436e4
62f2680c
300fa80f
204c0113
606c28d2
300f66d2
e80fe06c
00536006
03c36426
08040f56
0f36f016
80c3ff96
a56c41c3
228724cc
001129dc
740ca5c3
818c233c
333c2303
601c418c
611cffff
2683ff00
408c723c
37c37303
ffff341c
2b5413e4
b0dc13e4
c5a0000f
047370cf
05f2108c
6f20718c
03f3718f
2170218c
652029c3
043536e4
618f6720
34c302d3
20e44c6c
32c30354
4006ff93
43e44c6f
708f0354
40060073
29c3508f
d98068a0
0a4066bc
dd94c007
260b673c
60376006
208604c3
100c263c
0a3f38bc
336430e3
54dc6007
540c000c
818c323c
223c3203
001c418c
011cffff
3083ff00
32036832
542c740f
818c323c
223c3203
3083418c
32036832
544c742f
818c323c
223c3203
3083418c
32036832
546c744f
818c323c
223c3203
3083418c
32036832
548c746f
818c323c
223c3203
3083418c
408c133c
348f1203
2435c0a7
100c363c
75807f85
146c2c0f
fe7e033c
133c344c
542cfe7e
fe7e233c
740c23c3
ffff001c
b0ff011c
20063083
4500111c
323c31a3
a2c3fe7e
60a6516f
62126f20
6d0050cc
3ac370cf
b0ec2c8c
b6c3d4ac
22541be4
20542007
32c354cc
14ec3183
36e460c3
22e30694
318332c3
145432e4
12543fe7
211c4006
65008100
ffff601c
00ff611c
3be4b6c3
08c30735
debc25c3
00070a56
0ac33854
341c602c
60073fff
18c32454
12a4315c
35546007
f5244e24
1304315c
315c69d2
8c2f1324
702f6006
1327415c
68c300f3
1307465c
1327465c
323c702f
62d24004
083cf324
20461fc0
bebc4006
035309e0
41490ac3
6285716c
70cc716f
70cf7d85
14c308c3
0a0622bc
01330dd2
315c18c3
65d206a4
14c308c3
00933664
66bc04c3
01960a40
0f56f076
00000804
3f36f016
0077fd96
403781c3
2007c3c3
60076954
20066754
b8c32c0f
0004b21c
680c2bc3
103c08c3
6c80044e
28c390c3
6d00480c
103c08c3
6c80064e
433ca0c3
001c00f4
011c1074
3fe60000
09e2f6bc
106c301c
0000311c
6c0c6c0c
301c60b7
311c10a8
ac100000
c206e006
bfe617c3
0106343c
0b0d333c
7f5233c4
343c4383
0dc30347
0ae94180
2e540007
6f296097
17946007
6007692c
6b691494
11946007
06940067
21e448ec
64c30c35
29f20173
07940047
35e468ec
64c30434
007321c3
35c321c3
e207e025
80250554
53c312c3
c207fa13
001c0a94
011c1074
76bc0000
086609e4
64c306f3
0347463c
3dc30057
6cbc2e00
201c0a09
211c10a8
680c0000
000c08c3
680c0e61
1bc36e00
2c2f240c
6e00680c
000c09c3
680c0c4f
1ac36e00
2c6f240c
6e00680c
0eed00c6
6e00680c
2d8f2017
6e00680c
0d0f042c
6e00680c
640f1cc3
1074001c
0000011c
09e476bc
03960006
0f56fc76
00000804
0136f016
51c3ff96
4037454c
601700f3
03c38c2c
0a0ae8bc
40178037
3f5c59f2
774d0001
556f554f
0100053c
12c323c3
b0bc40c6
3f5c0891
76ed0001
576d23c3
63d2752c
4ccf4017
752f6006
10b0301c
0000311c
00268c0c
701c2006
711c10ac
63c30000
7c0c0293
680c4c80
692c6ed2
0a9435e4
680f6006
6c807c0c
4d2f4006
7fe5780c
9fe5780f
25050025
303c85d2
60e7fff0
0006e935
80760196
08040f56
0f36f016
42c3a0c3
41544007
680f6006
3d542007
e42c0410
a46cc44c
38847f00
133c6e80
301c00f4
311c10a8
2c100000
213c0006
39c30347
6ae94d00
1c546007
6007690c
6c4c1954
16943ae4
38e4680c
682c1394
109437e4
36e4684c
686c0d94
0a9435e4
001c500f
011c1074
76bc0000
000609e4
202501b3
0106313c
0b0d333c
7f5233c4
00251383
d4940207
f0760866
08040f56
0336f016
40c3fe96
72c381c3
400693c3
40cc440f
4007a246
416c5754
1f3c07c3
b12c0040
5abc4aa0
50c30a4e
4c940007
332c6057
60572f2f
4cef50ec
b10c6057
6057ad0f
2def31ec
69ec4057
1b9460c7
2a0f320c
522c6057
60574e2f
ae4fb24c
326c6057
60572e6f
4e8f528c
b2ac6057
6057aeaf
2ecf32cc
52ec6057
60574eef
af0fb30c
396c64c3
4ca0798c
40070057
9f5c1554
37c30007
0a0a6ebc
05d250c3
66bc0057
02130a40
c007d86c
0057ed94
20cc70cc
32e421c3
66bc0554
a2460a40
38c30073
05c30c0f
c0760296
08040f56
3f36f016
90c3ff96
72c3c1c3
df5ca3c3
408c0184
40374ed2
8f5c8006
18c30004
458c654c
91806d20
6037646c
00d377f2
654c19c3
8ca0258c
47e482c3
a0062f34
1fc30ac3
3dc34006
0a4e5abc
0ad260c3
a03700f3
05c3946c
0a4066bc
baf254c3
acd20893
4017748c
4c6f65d2
748f6017
548f00d3
346f2017
a0170053
4d4c6017
68a02d8c
47e49180
38c3dc14
ac6f63d2
19c30073
4006a46f
19c3548f
6f8064cc
648c64cf
603764d2
03935cc3
00079f5c
6017ff93
6d4c0d8c
47c36c20
023573e4
15c343c3
b0bc24c3
fe2008cb
4d8c6017
4d8f4a00
b600e7d2
6c6c6017
19c36037
e007648f
67c3e794
019606c3
0f56fc76
00000804
8e243016
604cf524
aaaa101c
aaaa111c
32e421c3
7fe72054
101c1e54
111cdddd
202fdddd
416c61ec
608720cc
323c0794
616f0140
fec0313c
323c00d3
616f0280
fd80313c
343c60cf
03c34004
f3246ad2
00f30006
4004343c
f32462d2
0a4066bc
08040c56
60090373
08946047
033c30c3
0812011e
02a34c29
60070293
00251154
03946027
01533fe5
323c4009
0180fff0
033521e4
00532006
20672520
0006e5b4
00000804
85961016
29b709f7
69374977
0f3c9f57
20060a30
0149201c
0891b0bc
04e12f5c
09dd2f5c
233c69d7
48f7420b
04612f5c
09e52f5c
233c69d7
48b7440b
04412f5c
09ed2f5c
783269d7
2f5c6877
2f5c0421
3f5c09f5
3f5c04a1
4957057d
420b323c
3f5c6837
3f5c0401
49570585
440b323c
3f5c67f7
3f5c03e1
4957058d
47b75832
03c13f5c
05953f5c
04812f5c
065d2f5c
233c6917
4777420b
03a12f5c
06652f5c
233c6917
4737440b
03812f5c
066d2f5c
78326917
2f5c66f7
2f5c0361
70090675
05bd3f5c
323c500c
66b7420b
03413f5c
05c53f5c
323c500c
6677440b
03213f5c
05cd3f5c
5832500c
3f5c4637
3f5c0301
500c05d5
608732c3
09d72894
2f3c302c
3f3c0d30
54bc0d70
00070a07
000ce4dc
85f7902c
02e12f5c
05dd2f5c
420b243c
2f5c45b7
2f5c02c1
243c05e5
4577440b
02a12f5c
05ed2f5c
783234c3
2f5c6537
2f5c0281
145305f5
3f5c7089
502c05dd
420b323c
3f5c64f7
3f5c0261
502c05e5
440b323c
3f5c64b7
3f5c0241
502c05ed
44775832
02213f5c
05f53f5c
2f5c5109
704c05fd
420b233c
2f5c4437
2f5c0201
704c0605
440b233c
2f5c43f7
2f5c01e1
704c060d
63b77832
01c12f5c
06152f5c
3f5c7189
506c061d
420b323c
3f5c6377
3f5c01a1
506c0625
440b323c
3f5c6337
3f5c0181
506c062d
42f75832
01613f5c
06353f5c
82b7908c
01412f5c
063d2f5c
420b243c
2f5c4277
2f5c0121
243c0645
4237440b
01012f5c
064d2f5c
783234c3
2f5c61f7
2f5c00e1
3f5c0655
3f5c04c1
49970f3d
420b323c
3f5c61b7
3f5c00c1
49970f45
440b323c
3f5c6177
3f5c00a1
49970f4d
41375832
00813f5c
0f553f5c
482c4997
3f5c40f7
3f5c0061
323c069d
60b7420b
00412f5c
06a52f5c
233c60d7
4077440b
00212f5c
06ad2f5c
783260d7
2f5c6037
2f5c0001
700606b5
0a1d3f5c
2f5c4006
2f5c0a25
2f5c0a2d
0f3c0a35
3f970a30
0a2096bc
08567b96
00000804
50c37016
64cc41c3
05b46267
66bc01c3
07130a40
139c301c
0000311c
6af26c0c
14c0303c
11b4201c
0000211c
23e4480c
4e242754
355cf524
6ed21c04
1c24355c
455c8c2f
60061c27
355c702f
60251c44
1c47355c
455c0133
455c1c07
702f1c27
655cc026
323c1c47
62d24004
053cf324
101c1fc0
40060080
09e0bebc
9ebc0073
0e560a26
00000804
0136f016
50c3f496
005c71c3
10c304c1
04c9055c
40ac303c
04d1155c
81ac313c
04d9255c
c1ac823c
64c39689
343c96a9
d6c9432c
81ac363c
403c16e9
18c3c1ac
06e4015c
02c01f3c
0b948087
60064706
0a4e5abc
54dc0007
62d70025
11f38def
60064706
0a4e5abc
b4dc0007
62d70024
8def80c6
655c42d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8a8f8c4c
655c42d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8aaf8c6c
655c42d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8acf8c8c
655c42d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8aef8cac
d70942d7
d72906c3
402c363c
303c1749
376981ac
c1ac313c
42d76a0f
64c39789
343c97a9
d7c9432c
81ac363c
303c17e9
6a2fc1ac
155c42d7
41c30101
0109155c
422c313c
0111455c
81ac343c
0119655c
c1ac363c
42d76a4f
0121055c
055c10c3
303c0129
155c40ac
313c0131
455c81ac
343c0139
6a6fc1ac
655c42d7
06c30181
0189655c
402c363c
0191055c
81ac303c
0199155c
c1ac313c
42d768ef
01a1455c
455c64c3
343c01a9
655c432c
363c01b1
055c81ac
303c01b9
690fc1ac
696c42d7
698f6285
228662d7
62d72ccf
7589cd6c
75a943c3
422c233c
0141455c
455c04c3
343c0149
055c402c
303c0151
155c81ac
313c0159
323cc1ac
780f81ac
255cf82f
42c30241
0249255c
422c323c
0251455c
81ac343c
0259055c
c1ac303c
155c784f
21c303c1
03c9155c
412c313c
03d1255c
81ac323c
03d9455c
c1ac343c
011c0006
30a35010
2006786f
255c388f
42c30241
0249255c
422c323c
0251455c
81ac343c
0259055c
c1ac103c
1f5c22b7
155c0141
42970265
420b323c
3f5c6277
355c0121
8297026d
440b043c
0f5c0237
055c0101
22970275
21f73832
00e12f5c
027d255c
03c1455c
455c04c3
343c03c9
055c402c
303c03d1
155c81ac
213c03d9
41b7c1ac
00c12f5c
03e5255c
433c6197
8177420b
00a14f5c
03ed455c
103c0197
2137440b
00811f5c
03f5155c
58324197
3f5c40f7
355c0061
301c03fd
311c1108
8c090000
0285455c
055c0c29
2c49028d
0295155c
255c4c69
580c029d
818c323c
223c3203
401c418c
411cffff
3483ff00
32036832
582c780f
818c323c
223c3203
3483418c
32036832
584c782f
818c323c
223c3203
3483418c
32036832
586c784f
818c323c
223c3203
3483418c
32036832
588c786f
818c323c
223c3203
3483418c
32036832
3689788f
36a921c3
412c313c
323c56c9
96e981ac
c1ac343c
13946087
0181155c
155c21c3
313c0189
255c412c
323c0191
455c81ac
343c0199
733cc1ac
02530140
0a21055c
055c10c3
303c0a29
155c40ac
313c0a31
255c81ac
323c0a39
733cc1ac
42d70080
353c88cc
60370180
20c602c3
37c324c3
0a3f38bc
233c30e3
323c800c
3203818c
418c223c
ffff401c
ff00411c
68323483
788f3203
06c3d689
363cd6a9
16c9402c
81ac303c
313c36e9
22d7c1ac
44946087
64c39709
343c9729
d749432c
81ac363c
203c1769
455cc1ac
64c304e1
04e9455c
432c343c
04f1655c
81ac363c
04f9055c
c1ac403c
0501655c
655c06c3
363c0509
055c402c
303c0511
655c81ac
363c0519
6037c1ac
011c0006
00770006
0521655c
655c06c3
363c0529
055c402c
303c0531
655c81ac
363c0539
60b7c1ac
34c308c3
0a22a0bc
055c0453
20c30a21
0a29055c
412c303c
0a31255c
81ac323c
0a39455c
c1ac343c
42d7670f
106c301c
0000311c
a8cc6c0c
665c68c3
c03731a4
08c38e4c
40c612c3
466435c3
80760c96
08040f56
f7963016
8e2410c3
036cf524
13540007
52c34009
323c4029
a04942ac
81ac353c
323c4069
501cc1ac
511c5020
25c35443
085432e4
4004343c
42dc6007
f324000d
301c1a33
311c139c
6c0c0000
6df261f7
11b4301c
0000311c
501c6c0c
511c12c0
25c30000
299432e4
243c674c
60074004
301c1f54
311cb50c
674f0014
04c1405c
405c54c3
343c04c9
505c42ac
353c04d1
105c81ac
013c04d9
42d2c1ac
021cf324
101c01fc
40061000
09e0bebc
40071373
000992dc
12d3f324
6007674c
0008f2dc
474f41d7
6237678c
129413e4
00e12f5c
0765205c
00e13f5c
076d305c
00e15f5c
0775505c
00e12f5c
077d205c
3f5c0433
305c0101
a2170765
420b253c
2f5c41b7
205c00c1
6217076d
440b533c
5f5ca177
505c00a1
42170775
41375832
00813f5c
077d305c
a7ac478c
67acabaf
205c4f8f
52c30781
0789205c
42ac323c
0791505c
81ac353c
0799205c
c1ac323c
fff0233c
3f5c40f7
305c0061
223c0785
40b7420b
00413f5c
078d305c
253ca0d7
4077440b
00212f5c
0795205c
783260d7
5f5c6037
505c0001
658c079d
28946187
0201505c
505c25c3
353c0209
205c412c
323c0211
505c81ac
353c0219
60a7c1ac
67060554
0427315c
a0260093
0427515c
1250201c
0000211c
6025680c
343c680f
62d24004
01c3f324
09f102bc
343c00b3
62d24004
0996f324
08040c56
f3967016
8e2410c3
036cf524
13540007
52c34009
323c4029
a04942ac
81ac353c
363cc069
201cc1ac
211c5020
52c35443
085435e4
4004343c
52dc6007
f3240012
301c2453
311c139c
6c0c0000
6df262f7
11b4301c
0000311c
601c6c0c
611c12c0
26c30000
299432e4
243c674c
60074004
301c1f54
311cb50c
674f0014
04c1405c
405c54c3
343c04c9
505c42ac
353c04d1
605c81ac
063c04d9
42d2c1ac
021cf324
101c01fc
40061000
09e0bebc
40071d93
000ea2dc
1cf3f324
6007674c
000e02dc
474f42d7
6337678c
129413e4
01616f5c
07a5605c
01612f5c
07ad205c
01613f5c
07b5305c
01615f5c
07bd505c
6f5c0433
605c0181
431707a5
420b323c
3f5c62b7
305c0141
a31707ad
440b653c
6f5cc277
605c0121
431707b5
42375832
01013f5c
07bd305c
a7ac478c
67acabaf
605c4f8f
26c307c1
07c9605c
412c363c
07d1205c
81ac323c
07d9505c
c1ac353c
fff0233c
3f5c41f7
305c00e1
623c07c5
c1b7420b
00c12f5c
07cd205c
533c61d7
a177440b
00a15f5c
07d5505c
d832c1d7
2f5cc137
205c0081
505c07dd
65c30221
0229505c
432c353c
0231605c
81ac363c
0239205c
c1ac323c
0140233c
accc67ec
60f76aa0
00616f5c
0225605c
420b333c
5f5c60b7
505c0041
c0d7022d
440b263c
2f5c4077
205c0021
60d70235
60377832
00015f5c
023d505c
6187658c
205c4a94
52c30201
0209205c
42ac323c
0211505c
81ac353c
0219605c
c1ac363c
035460a7
04d36706
05c1505c
505c65c3
353c05c9
605c432c
363c05d1
505c81ac
253c05d9
605cc1ac
56c305a1
05a9605c
42ac363c
05b1505c
81ac353c
05b9605c
c1ac363c
053423e4
215c4726
00930427
315c6926
201c0427
211c1250
680c0000
680f6025
4004343c
f32462d2
02bc01c3
00b309f1
4004343c
f32462d2
0e560d96
00000804
fa967016
f5242e24
4007436c
88091354
882954c3
42ac343c
353ca849
c86981ac
c1ac363c
5020401c
5443411c
35e454c3
313c0854
60074004
000d62dc
1a73f324
04c1625c
625c46c3
363c04c9
425c422c
343c04d1
525c81ac
453c04d9
301cc1ac
311c139c
6c0c0000
6df26177
11b4301c
0000311c
601c6c0c
611c12c0
56c30000
1a9435e4
213c634c
60074004
601c1054
611cb50c
c34f0014
f32442d2
1fc0043c
1000101c
bebc4006
13b309e0
b2dc4007
f3240009
634c1313
12dc6007
61570009
4f5c634f
425c00a1
5f5c07e5
525c00a1
6f5c07ed
625c00a1
3f5c07f5
325c00a1
4f5c07fd
425c00a1
5f5c0625
525c00a1
6f5c062d
625c00a1
3f5c0635
325c00a1
8909063d
892954c3
42ac343c
353ca949
c96981ac
c1ac463c
80078137
60261154
0205325c
00a14f5c
020d425c
00a15f5c
0215525c
00a16f5c
021d625c
60460793
0205325c
00814f5c
020d425c
00815f5c
0215525c
00816f5c
021d625c
0241425c
425c54c3
343c0249
525c42ac
353c0251
625c81ac
363c0259
533cc1ac
a0f7fff0
00616f5c
0245625c
420b453c
5f5c80b7
525c0041
c0d7024d
440b363c
3f5c6077
325c0021
80d70255
80379832
00015f5c
025d525c
6187618c
47061294
0427205c
1250201c
0000211c
6025680c
313c680f
62d24004
02bcf324
00b309f1
4004313c
f32462d2
0e560696
00000804
ff963016
8e2410c3
036cf524
13540007
52c34009
323c4029
a04942ac
81ac353c
323c4069
501cc1ac
511c5020
25c35443
075432e4
4004343c
6b546007
0d33f324
139c301c
0000311c
60376c0c
301c6df2
311c11b4
6c0c0000
12c0501c
0000511c
32e425c3
674c2894
4004243c
1f546007
b50c301c
0014311c
405c674f
54c304c1
04c9405c
42ac343c
04d1505c
81ac353c
04d9105c
c1ac013c
f32442d2
01fc021c
1000101c
bebc4006
067309e0
31544007
05f3f324
6007674c
40172854
3f5c474f
305c0001
5f5c0805
505c0001
2f5c080d
205c0001
3f5c0815
305c0001
658c081d
13946187
215c4826
201c0427
211c1250
680c0000
680f6025
4004343c
f32462d2
02bc01c3
00b309f1
4004343c
f32462d2
0c560196
00000804
40c33016
0201105c
105c21c3
313c0209
205c412c
323c0211
105c81ac
513c0219
4026c1ac
0205205c
305c6006
305c020d
305c0215
305c021d
305c0625
305c062d
305c0635
628d063d
62cd62ad
630d62ed
634d632d
638d636d
63cd63ad
305c63ed
305c0105
305c010d
305c0115
305c011d
305c0125
305c012d
305c0135
105c013d
21c305c1
05c9105c
412c313c
05d1205c
81ac323c
05d9105c
c1ac313c
e6bc63d2
245c0a4d
12c30541
0549245c
40ac323c
0551145c
81ac313c
0559245c
c1ac323c
04c367d2
0a13eebc
5abc0073
145c0a0f
21c30761
0769145c
412c313c
0771245c
81ac323c
0779145c
c1ac013c
ee940007
4ebc0073
245c0a10
12c307a1
07a9245c
40ac323c
07b1145c
81ac313c
07b9245c
c1ac023c
ee940007
07e1145c
145c21c3
313c07e9
245c412c
323c07f1
145c81ac
013c07f9
03d2c1ac
0a1194bc
0801245c
245c12c3
323c0809
145c40ac
313c0811
245c81ac
023c0819
03d2c1ac
0a128abc
1394a0a7
0941145c
145c21c3
313c0949
245c412c
323c0951
145c81ac
313c0959
63d2c1ac
366404c3
0901245c
245c12c3
323c0909
145c40ac
313c0911
245c81ac
323c0919
63d2c1ac
366404c3
08040c56
fc963016
105c50c3
21c30561
0569105c
412c313c
0571205c
81ac323c
0579105c
c1ac013c
255c4006
255c0565
255c056d
255c0575
255c057d
255c0585
255c058d
255c0595
06d3059d
301c804c
311caaaa
604faaaa
0a4066bc
0541155c
155c21c3
313c0549
255c412c
323c0551
155c81ac
313c0559
133cc1ac
20f7fff0
00612f5c
0545255c
420b113c
2f5c20b7
255c0041
60d7054d
440b133c
1f5c2077
155c0021
40d70555
40375832
00013f5c
055d355c
155c04c3
21c30541
0549155c
412c313c
0551255c
81ac323c
0559155c
c1ac313c
bb946007
0c560496
00000804
ff963016
4006646c
0010211c
60073283
000942dc
0221405c
405c54c3
343c0229
505c42ac
353c0231
205c81ac
423c0239
644cc1ac
7e9434e4
0241205c
205c52c3
323c0249
505c42ac
353c0251
505c81ac
253c0259
642cc1ac
6c9432e4
428d4006
42cd42ad
430d42ed
434d432d
438d436d
43cd43ad
205c43ed
205c0105
205c010d
205c0115
205c011d
205c0125
205c012d
205c0135
205c013d
205c0145
205c014d
205c0155
8109015d
812954c3
42ac343c
353ca149
216981ac
c1ac213c
4cd24037
205c4026
60060205
020d305c
0215305c
021d305c
80460213
0205405c
00015f5c
020d505c
00011f5c
0215105c
00012f5c
021d205c
305c6006
305c0625
305c062d
305c0635
405c063d
54c30801
0809405c
42ac343c
0811505c
81ac353c
0819105c
c1ac313c
021c6ad2
20060100
0a5738bc
14c30093
0a0cd6bc
0c560196
00000804
fc961016
005c40c3
10c302c1
02c9045c
40ac303c
02d1145c
81ac313c
02d9245c
c1ac323c
32dc6007
045c000b
10c302a1
02a9045c
40ac303c
02b1145c
81ac313c
02b9045c
c1ac203c
0241145c
145c01c3
313c0249
045c402c
303c0251
145c81ac
313c0259
23e4c1ac
000924dc
0a01145c
145c21c3
313c0a09
245c412c
323c0a11
045c81ac
303c0a19
6007c1ac
20061254
06c5145c
06cd145c
06d5145c
06dd145c
06e5145c
06ed145c
06f5145c
06fd145c
245c40c6
60060205
020d345c
0215345c
021d345c
0241045c
045c10c3
303c0249
145c40ac
313c0251
245c81ac
323c0259
133cc1ac
20f70010
00612f5c
0245245c
420b013c
1f5c00b7
145c0041
40d7024d
440b323c
3f5c6077
345c0021
00d70255
00371832
00011f5c
025d145c
5abc0073
245c0a0f
02c30761
0769245c
402c323c
0771045c
81ac303c
0779145c
c1ac013c
ee940007
0221245c
245c02c3
323c0229
045c402c
303c0231
04c381ac
0239245c
c1ac123c
0a0cd6bc
0941045c
045c10c3
303c0949
145c40ac
313c0951
245c81ac
323c0959
63d2c1ac
366404c3
08560496
00000804
ff963016
646c40c3
011c0006
30830010
42dc6007
245c000a
02c30221
0229245c
402c323c
0231045c
81ac303c
0239245c
c1ac523c
35e4644c
0008d4dc
0241245c
245c02c3
323c0249
045c402c
303c0251
045c81ac
203c0259
642cc1ac
7a9432e4
528d4006
52cd52ad
530d52ed
534d532d
538d536d
53cd53ad
245c53ed
245c0105
245c010d
245c0115
245c011d
245c0125
245c012d
245c0135
245c013d
245c0145
245c014d
245c0155
1109015d
112910c3
40ac303c
313c3149
516981ac
c1ac023c
0ad20037
345c6026
00060205
020d045c
0215045c
20460193
0205145c
00012f5c
020d245c
345c32c3
02c30215
021d045c
145c2006
145c0625
145c062d
145c0635
245c063d
02c30801
0809245c
402c323c
0811045c
81ac303c
0819145c
c1ac313c
043c66d2
20061000
0a5738bc
0901245c
245c02c3
323c0909
045c402c
303c0911
145c81ac
313c0919
68d2c1ac
366404c3
04c300b3
d6bc15c3
01960a0c
08040c56
0136f016
40c3f196
301c51c3
311c1110
6c0c0000
eebcec0c
60c309f8
346c6264
400601c3
0010211c
00070283
0011b2dc
0221245c
245c82c3
323c0229
245c442c
823c0231
345c81ac
233c0239
744cc42c
84dc32e4
31c30010
ffff341c
0ff4213c
0f5c4377
045c01a1
233c02e5
4337408c
01810f5c
02ed045c
145c2006
833c02f5
8f5cc08c
0f5c0167
045c0161
1f5c02fd
145c01a1
2f5c01e5
245c0181
600601ed
01f5345c
01fd045c
0161145c
145c21c3
313c0169
245c412c
323c0171
045c81ac
103c0179
01c3c1ac
1f5c22b7
145c0141
303c0305
6277420b
01213f5c
030d345c
440b103c
1f5c2237
145c0101
42970315
41f75832
00e13f5c
031d345c
045c00a6
20060205
020d145c
0215145c
021d145c
08e1245c
245c82c3
323c08e9
045c442c
303c08f1
145c81ac
313c08f9
63d2c1ac
366404c3
0a01245c
245c82c3
323c0a09
045c442c
303c0a11
145c81ac
313c0a19
6007c1ac
c0074554
375c1d54
36e405d9
363c1914
1c2c03c7
6d8b6c00
600763b7
1f5c1154
145c01c1
683206c5
2f5c61b7
245c00c1
600606cd
06d5345c
06dd345c
301c03d3
311c106c
6c0c0000
0ca96c0c
0cc910c3
40ac103c
217701c3
00a11f5c
06c5145c
483220c3
3f5c4137
345c0081
000606cd
06d5045c
06dd045c
145c2006
145c06e5
145c06ed
145c06f5
245c06fd
82c30241
0249245c
442c323c
0251045c
81ac303c
0259145c
c1ac213c
40f712c3
00612f5c
0265245c
420b813c
00478f5c
00410f5c
026d045c
440b213c
2f5c4077
245c0021
60d70275
60377832
00010f5c
027d045c
07e1145c
145c21c3
313c07e9
245c412c
323c07f1
045c81ac
303c07f9
6007c1ac
043c7e54
20060fc0
0a5738bc
31c30f13
211c4006
32830002
3d546007
0241045c
045c10c3
303c0249
145c40ac
313c0251
245c81ac
123c0259
045cc1ac
20c303c1
03c9045c
412c303c
03d1245c
81ac323c
03d9045c
c1ac303c
542c6c80
341431e4
041421e4
23e40673
245c3135
82c30221
0229245c
442c323c
0231045c
81ac303c
0239145c
c1ac313c
133c04c3
b0bcfff0
06b30a2c
33540007
0221245c
245c82c3
323c0229
045c442c
303c0231
145c81ac
213c0239
744cc1ac
215432e4
15c304c3
0a2096bc
21e40393
742ccf14
742f6025
15c304c3
0a2096bc
145c2026
40060205
020d245c
0215245c
021d245c
0625245c
062d245c
0635245c
063d245c
80760f96
08040f56
e296f016
51c340c3
1110301c
0000311c
ec0c6c0c
09f8eebc
626460c3
0006546c
0012011c
30c32083
a4dc23e4
045c0011
10c30221
0229045c
40ac303c
0231145c
81ac313c
0239045c
c1ac303c
13e4344c
001074dc
033c742c
07370010
03812f5c
0245245c
420b003c
2f5c06f7
245c0361
6717024d
440b033c
0f5c06b7
045c0341
47170255
46775832
03213f5c
025d345c
23c3746c
ffff241c
0ff4033c
3f5c0637
345c0301
023c02e5
05f7408c
02e13f5c
02ed345c
545ca006
323c02f5
65b7c08c
02c15f5c
02fd545c
03010f5c
01e5045c
02e12f5c
01ed245c
345c6006
545c01f5
345c01fd
345c0325
345c032d
345c0335
045c033d
20c30161
0169045c
412c303c
0171245c
81ac323c
0179545c
c1ac053c
057750c3
02a10f5c
0305045c
420b353c
3f5c6537
345c0281
053c030d
04f7440b
02610f5c
0315045c
58324557
3f5c44b7
345c0241
04c3031d
0a0cd6bc
545ca0a6
00060205
020d045c
0215045c
021d045c
0625045c
062d045c
0635045c
063d045c
08e1145c
145c21c3
313c08e9
245c412c
323c08f1
545c81ac
353c08f9
63d2c1ac
366404c3
0a01045c
045c10c3
303c0a09
145c40ac
313c0a11
245c81ac
323c0a19
6007c1ac
c0073d54
375c1554
36e405d9
363c1114
1c2c03c7
6d8b6c00
6ad26777
03a11f5c
06c5145c
64776832
02212f5c
301c02f3
311c106c
6c0c0000
aca96c0c
acc905c3
402c053c
043750c3
02010f5c
06c5045c
283215c3
2f5c23f7
245c01e1
600606cd
06d5345c
06dd345c
545ca006
545c06e5
545c06ed
545c06f5
045c06fd
10c307e1
07e9045c
40ac303c
07f1145c
81ac313c
07f9245c
c1ac323c
22dc6007
043c0010
20060fc0
0a5738bc
60061f73
0002311c
20e403c3
000ce4dc
233c742c
43b70010
01c13f5c
0245345c
420b123c
2f5c2377
245c01a1
6397024d
440b033c
0f5c0337
045c0181
23970255
22f73832
01612f5c
025d245c
23c3746c
ffff241c
0ff4033c
1f5c02b7
145c0141
523c02e5
a277408c
01210f5c
02ed045c
145c2006
523c02f5
a237c08c
01010f5c
02fd045c
01411f5c
01e5145c
01212f5c
01ed245c
345c6006
50c301f5
01fd545c
0161045c
045c10c3
303c0169
145c40ac
313c0171
245c81ac
523c0179
25c3c1ac
3f5ca1f7
345c00e1
053c0305
01b7420b
00c11f5c
030d145c
440b323c
3f5c6177
345c00a1
a1d70315
a137b832
00810f5c
031d045c
145c2006
145c0325
145c032d
145c0335
245c033d
52c30221
0229245c
42ac323c
0231545c
81ac353c
0239045c
c1ac303c
0010233c
3f5c40f7
345c0061
023c0225
00b7420b
00411f5c
022d145c
440b323c
5f5c6077
545c0021
00d70235
00371832
00011f5c
023d145c
245c4086
60060205
020d345c
0215345c
021d345c
0625345c
062d345c
0635345c
063d345c
0221545c
545c05c3
353c0229
045c402c
303c0231
126481ac
c1ac313c
133c04c3
b0bcfff0
05130a2c
31c3346c
211c4006
32830010
20546007
0221045c
045c20c3
303c0229
245c412c
323c0231
045c81ac
203c0239
744cc1ac
0e5432e4
400631c3
0002211c
64d23283
6025742c
04c3742f
96bc15c3
1e960a20
08040f56
0136f016
60c3de96
04c1005c
065c10c3
303c04c9
165c40ac
313c04d1
265c81ac
823c04d9
065cc1ac
10c307a1
07a9065c
40ac303c
07b1165c
81ac313c
07b9265c
c1ac123c
62dc2007
e7ec002e
0301065c
065c10c3
303c0309
165c40ac
213c0311
065c81ac
10c302e1
02e9065c
40ac303c
02f1165c
81ac313c
02f9065c
c1ac303c
0319165c
c12c213c
023523e4
165c23c3
01c30321
0329165c
402c313c
0331065c
81ac303c
0339165c
c1ac313c
23e42006
29a00235
7d857ccc
c0dc13e4
065c002a
10c305c1
05c9065c
40ac303c
05d1165c
81ac313c
05d9065c
c1ac203c
05a1165c
165c01c3
313c05a9
065c402c
303c05b1
165c81ac
313c05b9
23e4c1ac
0028b1dc
0981165c
165c21c3
313c0989
265c412c
323c0991
065c81ac
303c0999
63d2c1ac
366406c3
05e1165c
165c21c3
313c05e9
265c412c
323c05f1
065c81ac
103c05f9
2877c1ac
0ff4273c
073c41b7
0177408c
808c273c
073c4137
00f7c08c
20072857
265c2254
02c30601
0609265c
402c323c
0611065c
81ac303c
0619165c
c1ac313c
2f5cec4f
265c00c1
3f5c0605
365c00a1
0f5c060d
065c0081
1f5c0615
165c0061
0bd3061d
00c12f5c
05e5265c
03c36157
00ff041c
1f5c0837
165c0401
411705ed
341c32c3
67f700ff
03e10f5c
05f5065c
00611f5c
05fd165c
00c12f5c
0605265c
04013f5c
060d365c
0615065c
061d165c
0641265c
265c02c3
323c0649
065c402c
303c0651
165c81ac
213c0659
12c3c1ac
2f5c47b7
265c03c1
013c0625
0777420b
03a10f5c
062d065c
440b213c
2f5c4737
265c0381
67970635
66f77832
03610f5c
063d065c
04211f5c
0665165c
265c21c3
31c3066d
0675365c
065c01c3
101c067d
111ceeee
3c4feeee
05c1265c
265c02c3
323c05c9
065c402c
303c05d1
165c81ac
313c05d9
033cc1ac
06b70010
03411f5c
05c5165c
420b303c
0f5c6677
065c0321
269705cd
440b213c
2f5c4637
265c0301
669705d5
65f77832
02e10f5c
05dd065c
0321165c
165c21c3
313c0329
265c412c
323c0331
065c81ac
303c0339
3cccc1ac
033c6c80
05b7fec0
02c11f5c
0325165c
420b303c
0f5c6577
065c02a1
2597032d
440b213c
2f5c4537
265c0281
65970335
64f77832
02610f5c
033d065c
0401165c
165c21c3
313c0409
265c412c
323c0411
065c81ac
303c0419
233cc1ac
44b70010
02413f5c
0405365c
420b123c
2f5c2477
265c0221
6497040d
440b033c
0f5c0437
065c0201
24970415
23f73832
01e12f5c
041d265c
0421065c
065c10c3
303c0429
165c40ac
313c0431
265c81ac
323c0439
1cccc1ac
233c6c00
43b7fec0
01c13f5c
0425365c
420b123c
2f5c2377
265c01a1
6397042d
440b033c
0f5c0337
065c0181
23970435
22f73832
01612f5c
043d265c
10c31a89
303c1aa9
3ac940ac
81ac313c
323c5ae9
6087c1ac
7def4694
21c33b09
313c3b29
5b49412c
81ac323c
203c1b69
165cc1ac
01c304e1
04e9165c
402c313c
04f1065c
81ac303c
04f9165c
c1ac413c
0501065c
065c10c3
303c0509
165c40ac
313c0511
065c81ac
303c0519
6037c1ac
111c2006
20770006
0521065c
065c10c3
303c0529
165c40ac
313c0531
065c81ac
303c0539
60b7c1ac
17c308c3
a0bc34c3
13f30a22
3def20c6
0a21265c
265c02c3
323c0a29
065c402c
303c0a31
165c81ac
313c0a39
4c4cc1ac
065c5e8f
10c30a21
0a29065c
40ac303c
0a31165c
81ac313c
0a39265c
c1ac323c
1eaf0c6c
0a21165c
165c21c3
313c0a29
265c412c
323c0a31
065c81ac
303c0a39
2c8cc1ac
265c3ecf
02c30a21
0a29265c
402c323c
0a31065c
81ac303c
0a39165c
c1ac313c
5eef4cac
10c31b09
303c1b29
3b4940ac
81ac313c
323c5b69
7e0fc1ac
10c31b89
303c1ba9
3bc940ac
81ac313c
323c5be9
7e2fc1ac
0101065c
065c10c3
303c0109
165c40ac
313c0111
265c81ac
323c0119
7e4fc1ac
0121065c
065c10c3
303c0129
165c40ac
313c0131
265c81ac
323c0139
7e6fc1ac
0a21065c
065c10c3
303c0a29
165c40ac
313c0a31
265c81ac
323c0a39
7f0fc1ac
106c301c
0000311c
bccc6c0c
005c08c3
003731a4
08c38e4c
40c617c3
466435c3
07c1165c
165c21c3
313c07c9
265c412c
323c07d1
065c81ac
303c07d9
233cc1ac
42b7fff0
01413f5c
07c5365c
420b123c
2f5c2277
265c0121
629707cd
440b033c
0f5c0237
065c0101
229707d5
21f73832
00e12f5c
07dd265c
0f40063c
38bc2006
22960a57
0f568076
00000804
0336f016
70c3da96
256c51c3
323c440c
3203818c
418c223c
ffff001c
ff00011c
033c3083
0203408c
442c040f
818c323c
223c3203
401c418c
411cffff
3483ff00
32036832
233c642f
74cc808c
80dc32e4
80c30011
ffff841c
408c383c
933c3884
301c00f4
311c11b4
6c0c0000
301c6cd2
311c139c
6c0c0000
073c66f2
3fe60e00
09e2f6bc
0b60393c
3a1d673c
c00746c3
75ec3394
1b9460c7
15e4375c
17546007
6ccc772c
011c0006
3083ff00
32e420c3
301c0e54
311c106c
6c0c0000
07c38e2c
400615c3
0104211c
466436c3
11b4301c
0000311c
60076c0c
000d32dc
139c301c
0000311c
60076c0c
000cb4dc
0e00073c
09e476bc
110918b3
112910c3
40ac303c
313c3149
516981ac
c1ac323c
289438e4
21c33389
313c33a9
53c9412c
81ac323c
303c13e9
34ccc1ac
033c6c80
08f7ff80
04611f5c
303c338d
68b7420b
04410f5c
28d713ad
440b213c
2f5c4877
53cd0421
783268d7
0f5c6837
13ed0401
145c0253
21c30261
0269145c
412c313c
0271245c
81ac323c
0279045c
c1ac403c
bc9446e4
11b4301c
0000311c
6bd26c0c
139c301c
0000311c
65f26c0c
0e00073c
09e476bc
02c35109
323c5129
1149402c
81ac303c
313c3169
38e4c1ac
75ec1f54
609460c7
15e4375c
5c546007
6ccc772c
011c0006
3083ff00
32e420c3
301c5354
311c106c
6c0c0000
07c38e2c
400615c3
0104211c
46646006
2e2408b3
1009f524
102920c3
412c303c
323c5049
106981ac
c1ac303c
5020201c
5544211c
30e402c3
245c3554
72c30121
0129245c
43ac323c
0131745c
81ac373c
0139045c
c1ac303c
0010733c
0f5ce7f7
045c03e1
373c0125
67b7420b
03c17f5c
012d745c
203c07d7
4777440b
03a12f5c
0135245c
783267d7
7f5c6737
745c0381
313c013d
62d24004
05c3f324
0a4066bc
045c3e93
20c30381
0389045c
412c303c
0391245c
81ac323c
0399045c
c1ac603c
0b60293c
2a1d373c
40e403c3
375c0654
63f20744
2b9d473c
02c1245c
245c72c3
323c02c9
745c43ac
373c02d1
245c81ac
023c02d9
0007c1ac
638c7054
03e46937
40060b94
02c5245c
02cd245c
02d5245c
02dd245c
3f5c0433
345c0481
e91702c5
420b273c
2f5c46f7
245c0361
691702cd
440b733c
7f5ce6b7
745c0341
491702d5
46775832
03213f5c
02dd345c
e3ac438c
63acebaf
245c4f8f
72c302e1
02e9245c
43ac323c
02f1745c
81ac373c
02f9245c
c1ac323c
fff0233c
3f5c4637
345c0301
223c02e5
45f7420b
02e13f5c
02ed345c
273ce617
45b7440b
02c12f5c
02f5245c
78326617
7f5c6577
745c02a1
400602fd
201c434f
211c1250
680c0000
680f6025
ac0f63ec
4004313c
f32462d2
305c6006
02bc0427
2ad309f1
0221745c
745c27c3
373c0229
245c412c
323c0231
745c81ac
373c0239
753cc1ac
e0f70ff4
408c753c
753ce0b7
e077808c
c08c753c
6007e037
000df2dc
0241245c
245c72c3
323c0249
745c43ac
373c0251
245c81ac
323c0259
ac2fc1ac
00613f5c
0245345c
00417f5c
024d745c
00212f5c
0255245c
00013f5c
025d345c
545c142f
75c301e1
01e9545c
43ac353c
01f1745c
81ac373c
01f9045c
c1ac303c
0010533c
7f5ca977
745c04a1
253c01e5
4537420b
02813f5c
01ed345c
440b753c
0f5ce4f7
045c0261
495701f5
44b75832
02413f5c
01fd345c
0201545c
545c75c3
353c0209
745c43ac
373c0211
045c81ac
303c0219
213cc1ac
29574004
53e451c3
745c7935
07c30221
0229745c
402c373c
0231045c
81ac303c
0239145c
c1ac013c
345c6089
a0a90225
022d545c
745ce0c9
20e90235
023d145c
01e1545c
545c75c3
353c01e9
745c43ac
373c01f1
145c81ac
313c01f9
733cc1ac
e477fff0
02211f5c
01e5145c
420b573c
7f5ca437
745c0201
245701ed
440b313c
3f5c63f7
345c01e1
a45701f5
a3b7b832
01c17f5c
01fd745c
0121145c
145c51c3
313c0129
545c42ac
353c0131
745c81ac
373c0139
533cc1ac
a3770010
01a17f5c
0125745c
420b353c
5f5c6337
545c0181
e357012d
440b173c
1f5c22f7
145c0161
63570135
62b77832
01415f5c
013d545c
f32442d2
0a4066bc
40070bf3
f3245d54
7f5c0b73
745c0061
00970225
241c20c3
427700ff
01217f5c
022d745c
20c30057
00ff241c
7f5c4237
745c0101
0f5c0235
045c0001
2f5c023d
245c0061
7f5c0245
745c0121
0f5c024d
045c0101
2f5c0255
245c0001
742f025d
01e1545c
545c75c3
353c01e9
745c43ac
373c01f1
045c81ac
303c01f9
533cc1ac
a1f70010
00e17f5c
01e5745c
420b253c
3f5c41b7
345c00c1
753c01ed
e177440b
00a10f5c
01f5045c
583241d7
3f5c4137
345c0081
313c01fd
62d24004
c3d2f324
666404c3
c0762696
08040f56
0136f016
50c3fc96
005c71c3
10c304c1
04c9055c
40ac303c
04d1155c
81ac313c
04d9255c
c1ac823c
64c39689
343c96a9
d6c9432c
81ac363c
403c16e9
18c3c1ac
06e4015c
00c01f3c
0b948087
60064706
0a4e5abc
b4dc0007
60d7001d
11f38def
60064706
0a4e5abc
14dc0007
60d7001d
8def80c6
655c40d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8a8f8c4c
655c40d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8aaf8c6c
655c40d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8acf8c8c
655c40d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8aef8cac
d70940d7
d72906c3
402c363c
303c1749
376981ac
c1ac313c
40d76a0f
64c39789
343c97a9
d7c9432c
81ac363c
303c17e9
6a2fc1ac
155c40d7
41c30101
0109155c
422c313c
0111455c
81ac343c
0119655c
c1ac363c
40d76a4f
0121055c
055c10c3
303c0129
155c40ac
313c0131
455c81ac
343c0139
6a6fc1ac
655c40d7
06c30181
0189655c
402c363c
0191055c
81ac303c
0199155c
c1ac313c
40d768ef
01a1455c
455c64c3
343c01a9
655c432c
363c01b1
055c81ac
303c01b9
690fc1ac
696c40d7
698f6285
228660d7
60d72ccf
7589cd6c
75a943c3
422c233c
0141455c
455c04c3
343c0149
055c402c
303c0151
155c81ac
313c0159
323cc1ac
780f81ac
40067c6c
0010211c
62d23283
782f7c4c
184f1c2c
03c1455c
455c14c3
343c03c9
155c40ac
313c03d1
255c81ac
123c03d9
6006c1ac
5014311c
580c13a3
818c323c
223c3203
401c418c
411cffff
3483ff00
32036832
582c780f
818c323c
223c3203
3483418c
32036832
303c782f
3003818c
418c203c
68323483
784f3203
818c313c
213c3103
3483418c
32036832
4006786f
9689588f
96a904c3
402c343c
303c16c9
36e981ac
c1ac313c
13946087
0181455c
455c04c3
343c0189
055c402c
303c0191
155c81ac
313c0199
733cc1ac
02530140
0a21255c
255c42c3
323c0a29
455c422c
343c0a31
055c81ac
303c0a39
733cc1ac
40d70080
353c88cc
60370180
20c602c3
37c324c3
0a3f38bc
233c30e3
323c800c
3203818c
418c223c
ffff101c
ff00111c
68323183
788f3203
42c35689
323c56a9
96c9422c
81ac343c
363cd6e9
20d7c1ac
44946087
42c35709
323c5729
9749422c
81ac343c
263cd769
055cc1ac
40c304e1
04e9055c
422c303c
04f1455c
81ac343c
04f9655c
c1ac463c
0501055c
055c60c3
303c0509
655c432c
363c0511
055c81ac
303c0519
6037c1ac
311c6006
60770006
0521655c
655c06c3
363c0529
055c402c
303c0531
655c81ac
363c0539
60b7c1ac
34c308c3
0a22a0bc
055c0453
20c30a21
0a29055c
412c303c
0a31255c
81ac323c
0a39455c
c1ac343c
40d7670f
106c301c
0000311c
a8cc6c0c
665c68c3
c03731a4
08c38e4c
40c612c3
466435c3
80760496
08040f56
0736f016
70c3f396
62c341c3
af5c23c3
64ec02e4
650c63d2
716c68f2
716f7d85
628570cc
447370cf
533c656c
a56ffec0
628564cc
052c64cf
51e410c3
002180dc
ffff341c
011c0006
30a34500
740f32a3
06c4275c
852c323c
323c742f
375c0010
459706c7
133c6557
344fc12c
0cac70ec
323c540c
3203818c
418c823c
ffff201c
ff00211c
68323283
740f3803
323c542c
3203818c
418c823c
ffff201c
ff00211c
68323283
742f3803
818c313c
213c3103
101c418c
111cffff
3183ff00
32036832
303c744f
3003818c
418c203c
68323183
746f3203
818c363c
263c3603
3183418c
32036832
4006748f
04c34037
42862086
38bc6006
30e30a3f
236423c3
818c323c
223c3203
001c418c
011cffff
3083ff00
32036832
31a3344c
30ec744f
400744a9
001752dc
04f004cc
508356c3
0b9458e4
36c320e3
32e43283
44ac0654
63e432c3
000814dc
0854dfe7
129458e4
36c320e3
32e43283
e2b70d94
01370086
101c8237
111cffff
21b70000
41f75fe6
175c11b3
21c325e4
b2dc62e4
a0060017
8100511c
001c7a80
011cffff
10c300ff
d9dc31e4
36c30014
211c4006
3283f000
511ca006
95c3e000
4a9439e4
0100001c
36c301b7
ffff101c
007f111c
40063183
5e00211c
61f732a3
106c301c
0000311c
6c0c6c0c
40062de9
375c0113
333c13e4
36e42a1d
40250554
f81421e4
375c0273
333c1464
6ed22a1d
1f3c04c3
275c0300
600606e4
0a0a06bc
07c305f2
18bc2317
e2b70a07
01370006
50ec8237
70cc42f7
51c3292c
c9dc35e4
175c0009
20071284
001202dc
4000a31c
001184dc
dc4c2353
72dcc007
363c0011
6f00408c
01f4933c
80c30e24
393cf524
273c0f30
40073a1d
690c4754
449436e4
31c3292c
35a3a94c
15546007
094c21b7
383c01f7
62d24004
e2b7f324
21372006
50ec8237
70cc42f7
95c3a92c
35dc39e4
0c53000e
345c702f
2d69fbc4
20f72272
00615f5c
698cad6d
6bf2a026
303c898f
60074004
000e82dc
1cb3f324
31c3a025
3df22c2c
01c38c2f
00c7531c
098c0535
698f602c
383c202f
62d24004
0007f324
000c54dc
383c1a13
12c34004
f3246bd2
011312c3
36e4650c
24ac0754
e2dc12e4
39f2000b
652c1773
454c03c3
000702a3
61b72554
61f7654c
f5246e24
0f30293c
2b9d173c
0400341c
f32462d2
a006e2b7
8237a137
42f750ec
092c70cc
31e410c3
175c0b35
20071284
000902dc
4000a31c
000884dc
6a0c1153
ce2411b3
345cf524
ad69fbc4
a0b7a272
00412f5c
102f4d6d
a026658c
858f6bf2
4004363c
32dc6007
f3240008
a0251013
4c2c32c3
8c2f5df2
531c02c3
053500c7
a02c058c
402fa58f
4004363c
f32462d2
60940007
893c0d93
383c0f30
07c3100c
56643d80
55940007
373c18c3
4ccc1a1d
092fc90f
301c094f
311c106c
6c0c0000
6d496c0c
084f682f
696f70ec
345c102f
ad69fbc4
a077a272
00210f5c
898f0d6d
2364375c
16c307c3
366450ec
a0060813
8100511c
001c7a80
011cffff
50c300ff
053535e4
30c304ac
109463e4
1f3c04c3
275c0300
600606e4
0a0a06bc
19940007
231707c3
0a0718bc
e2b70293
82374137
70cc22f7
95c3a52c
0f3539e4
1284175c
a31c28d2
05544000
01000f3c
01f31664
e8bc04c3
01730a0a
0f3c660c
36640100
575c00d3
a0072304
fe739794
e0760d96
08040f56
3f36f016
40c3ef96
0e00a03c
3fe60ac3
09e2f6bc
045c0026
64c308a7
0000801c
00c09f3c
106cc01c
0000c11c
02c0bf3c
2561165c
4e542007
2744365c
4a546007
42668277
383c40f7
321c0447
f18004a8
365ce2b7
09c32744
82773664
60f76026
2744365c
366409c3
00468277
365c00f7
09c32744
565c3664
02f32644
111c2006
22f7ff02
43374006
63776026
000674ac
ff00011c
63b730a3
640c1cc3
04c36e6c
27c31bc3
b4cc3664
e994a007
3144345c
10546007
211c4006
42f7ff02
a377a337
63b76026
600c0cc3
04c36e6c
27c31bc3
821c3664
c8850001
0002831c
b43caa94
df3c1fc0
6e240400
4004933c
03c0cf3c
00c08f3c
106c701c
0000711c
76bc0ac3
5fe609e4
0bc34037
402612c3
2abc3dc3
0ac309e0
f6bc3fe6
641709e2
0008341c
02d36ff2
642cf524
0927345c
345c63f2
39c30947
f32462d2
3abc04c3
145c0a07
31f20924
63926417
60076437
3f5cd854
67320201
345c6ad2
04c31be4
64173664
64376792
cb546007
341c6417
60070100
345c2854
600715e4
145c1554
28d22644
60676788
7c0c0594
04c36e8c
145c3664
28d22864
60676788
7c0c0594
04c36e8c
345c3664
63d21624
366404c3
1bc4345c
04c363d2
64173664
64376892
9f546007
341c6417
60070001
345c3b54
63d22324
366404c3
2444345c
04c363d2
345c3664
63d212c4
366404c3
14c4345c
04c363d2
345c3664
63d21ba4
366404c3
15e4345c
7c0c66d2
04c36e8c
36642006
1644345c
04c363d2
345c3664
65d215e4
6eac7c0c
366404c3
15e4345c
7c0c65d2
04c36ecc
64173664
64376092
12dc6007
6417fff6
0010341c
345c66d2
63d22344
366404c3
341c6417
66d20020
2464345c
04c363d2
64173664
0002341c
345c65d2
04c312a4
64173664
0004341c
345c65d2
04c315a4
64173664
0040341c
345c65d2
04c314e4
64173664
0400341c
2b546007
2561345c
12546007
01068277
101c00f7
21770100
211c4026
41b75e00
4a80343c
345c62b7
08c32744
345c3664
60072781
82771254
00f70106
0100101c
40262177
5e00211c
343c41b7
62b74ec0
2964345c
366408c3
341c6417
64c30800
6007a006
05131294
62468277
353c60f7
321c0447
718004a8
cf5c62b7
365c0107
08c32524
a0253664
2561065c
0b0d303c
233c33c4
4077f88c
00213f5c
600623c3
02d4a027
02c36026
00b70383
00413f5c
6007c885
6417da94
1000341c
32dc6007
345cffed
04c32524
d9b33664
fc761196
08040f56
3f36f016
b0c3c096
65ec71c3
6087472c
523c0994
a23c00c0
201c0100
4eb70218
523c0133
a23c0080
801c0180
8f5c04c4
7ccc0747
0007af5c
20c607c3
35c323c3
0a3f38bc
336430e3
14dc6007
3d70005e
400c09c3
818c323c
223c3203
101c418c
111cffff
3183ff00
32036832
402c600f
818c323c
223c3203
3183418c
32036832
404c602f
818c323c
223c3203
3183418c
32036832
406c604f
818c323c
223c3203
3183418c
408c133c
206f1203
323c408c
3203818c
418c223c
ffff001c
ff00011c
68323083
29c33203
313c688f
133ce08c
2007ffb0
7d6c1354
0140033c
1abc2212
0eb70a0b
7dec0bf2
0218101c
60872eb7
801c0554
8f5c04c4
09c30747
c3c3600c
ffffc41c
808c833c
07278f5c
408c3c3c
d33c3c84
3d3c00f4
0bc30ca0
3a1d803c
200718c3
000ec2dc
418908c3
41a912c3
40ac323c
313c21c9
41e981ac
c1ac323c
94dc3ce4
205c000c
12c30141
0149205c
40ac323c
0151105c
81ac313c
0159205c
c1ac323c
21c32e57
54dc32e4
2289000b
22a921c3
412c313c
323c42c9
22e981ac
c1ac213c
13c37dec
54dc21e4
2309000a
60b76329
c3698349
0e944087
323c4097
343c40ac
363c81ac
340cc1ac
32e421c3
000924dc
40970853
40ac323c
81ac343c
c1ac363c
21c3340c
54dc32e4
23890008
23a921c3
412c313c
323c43c9
23e981ac
c1ac313c
12c3542c
759431e4
0101205c
205c12c3
323c0109
105c40ac
313c0111
205c81ac
323c0119
344cc1ac
32e421c3
105c6294
21c30121
0129105c
412c313c
0131205c
81ac323c
0139105c
c1ac313c
12c3546c
4f9431e4
0ca03d3c
023c2bc3
19c33b9d
4006646c
0002211c
60073283
3f5c3d54
305c0741
2e970165
420b213c
2f5c4df7
205c06e1
6e97016d
440b833c
06c78f5c
06c11f5c
0175105c
58324e97
3f5c4d77
305c06a1
2e97017d
128d213c
2f5c4d37
205c0681
6d1701c5
420b833c
06678f5c
06611f5c
01cd105c
323c4d17
6cb7440b
06413f5c
01d5305c
38322d17
2f5c2c77
205c0621
17c301dd
0a2f84bc
0004a59c
0701105c
105c21c3
313c0709
205c412c
323c0711
105c81ac
013c0719
04d2c1ac
a4dc08e4
80c3fff1
606c09c3
111c2006
31830012
211c4006
02c30002
069430e4
315c1bc3
60071ca4
29c31094
0006686c
0004011c
60073083
0042f2dc
315c1bc3
60071ca4
004292dc
2ac3740c
10c3080c
159431e4
082c742c
31e410c3
744c1094
10c3084c
0b9431e4
086c746c
31e410c3
4e570694
3ce432c3
004502dc
205c0bc3
62c31ca4
3ce4780c
004034dc
106c301c
0000311c
6c0c6c0c
40074f49
301c1454
311c1110
4c0c0000
6f0b680c
0b9460a7
0884325c
17c3184c
30c33664
60073264
0042c2dc
8007984c
003442dc
606c09c3
111c2006
31830004
b4dc6007
7dec0033
0201145c
0209245c
0211045c
0219845c
25946087
40ac323c
81ac303c
c1ac383c
35946087
31c3340c
211c4006
3283e000
32dc32e4
7cec0040
0cec4ccc
328331c3
079430e4
31c322e3
32e43283
003f62dc
32dc10e4
3fe7003f
7df31a94
40ac323c
81ac303c
c1ac383c
11946087
106c301c
0000311c
6eec6c0c
366405c3
000630c3
4000011c
31e410c3
003d82dc
08c1245c
245c82c3
323c08c9
045c442c
303c08d1
145c81ac
313c08d9
67d2c1ac
17c304c3
00273664
003c24dc
784f6006
60877dec
1f894c94
0185045c
145c3fa9
5fc9018d
0195245c
345c7fe9
0bc3019d
243c340c
343c0300
54bc0340
0dd20a07
045c1409
342901a5
01ad145c
245c5449
746901b5
01bd345c
128d0086
32ad2006
32ed32cd
530d5409
732d7429
134d1449
336d3469
6d2c7cec
fd80833c
06078f5c
06010f5c
283c120d
4bf7420b
05e13f5c
183c722d
2bb7440b
05c12f5c
38c3524d
6b777832
05a10f5c
0cd3126d
328d20c6
52ad4006
52ed52cd
730d7409
132d1429
334d3449
536d5469
738d7489
13ad14a9
33cd34c9
53ed54e9
345c7509
15290105
010d045c
145c3549
55690115
011d245c
345c7589
15a90125
012d045c
145c35c9
55e90135
013d245c
6d2c7cec
fc40133c
2f5c2b37
520d0581
420b813c
05678f5c
05610f5c
213c122d
4ab7440b
05413f5c
0b17724d
0a771832
05211f5c
275c326d
245c0301
375c0a25
345c0309
075c0a2d
045c0311
175c0a35
145c0319
5f890a3d
0185245c
345c7fa9
1fc9018d
0195045c
145c3fe9
2f5c019d
245c0721
6e570145
6a376832
05010f5c
014d045c
145c2006
145c0155
29c3015d
245c4889
39c30245
345c6ca9
09c3024d
045c00c9
19c30255
145c24e9
4e97025d
341c32c3
69f700ff
04e10f5c
0165045c
213c2e97
49b7420b
04c12f5c
016d245c
833c6e97
8f5c440b
0f5c04a7
045c04a1
2e970175
29373832
04812f5c
017d245c
833c6e97
8f5c328d
0f5c0467
045c0461
283c01c5
48b7420b
04413f5c
01cd345c
440b183c
2f5c2877
245c0421
38c301d5
68377832
04010f5c
01dd045c
02e1145c
145c21c3
313c02e9
245c412c
323c02f1
045c81ac
103c02f9
27f7c1ac
03e11f5c
01e5145c
323c47d7
67b7420b
03c13f5c
01ed345c
103c07d7
2777440b
03a11f5c
01f5145c
583247d7
3f5c4737
345c0381
0f5c01fd
045c04e1
1f5c0305
145c04c1
2f5c030d
245c04a1
3f5c0315
345c0481
0006031d
0325045c
032d045c
0335045c
033d045c
0ca01d3c
223c2bc3
4e371a1d
0ff4843c
00878f5c
408c043c
808c543c
c08c343c
4e1760f7
92dc4007
3f5c0008
345c0701
323c0705
66f7420b
03612f5c
070d245c
833c6e17
8f5c440b
2f5c0347
245c0341
6e170715
66777832
03212f5c
071d245c
323c2bc3
235c1a1d
82c30721
0729235c
442c923c
0731235c
84ac923c
0739235c
c4ac823c
03078f5c
03013f5c
0725345c
420b383c
2f5c65f7
245c02e1
883c072d
8f5c440b
2f5c02c7
245c02c1
66170735
65777832
02a12f5c
073d245c
323c2bc3
235c1a1d
82c30721
0729235c
442c923c
0731235c
84ac823c
0739235c
c42c323c
00812f5c
0705235c
0ff4803c
02878f5c
02810f5c
070d035c
0ff4853c
02678f5c
02610f5c
0715035c
00612f5c
071d235c
303c0bc3
1f5c1a1d
135c0081
2f5c0725
235c0281
0f5c072d
035c0261
1f5c0735
135c0061
0573073d
00812f5c
0705245c
0ff4803c
02478f5c
02410f5c
070d045c
0ff4353c
0f5c6477
045c0221
2f5c0715
245c0061
3f5c071d
345c0081
0f5c0725
045c0241
2f5c072d
245c0221
3f5c0735
345c0061
0bc3073d
1b9d403c
07c3b82c
0a4066bc
0201145c
145c21c3
313c0209
245c412c
323c0211
045c81ac
303c0219
6087c1ac
000a34dc
0241245c
245c82c3
323c0249
045c442c
303c0251
145c81ac
313c0259
833cc1ac
8f5c0010
0f5c0207
045c0201
283c0245
43f7420b
01e13f5c
024d345c
440b183c
2f5c23b7
245c01c1
38c30255
63777832
01a10f5c
025d045c
0221145c
145c21c3
313c0229
245c412c
323c0231
045c81ac
303c0239
233cc1ac
43370010
01813f5c
0225345c
420b123c
2f5c22f7
245c0161
6317022d
440b833c
01478f5c
01410f5c
0235045c
38322317
2f5c2277
245c0121
045c023d
10c30641
0649045c
40ac303c
0651145c
81ac313c
0659245c
c1ac823c
01078f5c
01013f5c
0625345c
420b183c
2f5c21f7
245c00e1
883c062d
8f5c440b
0f5c00c7
045c00c1
22170635
21773832
00a12f5c
063d245c
345c6006
345c0665
345c066d
345c0675
045c067d
10c30221
0229045c
40ac303c
0231145c
81ac313c
0239245c
c1ac323c
133c04c3
b0bcfff0
a0070a2c
000f12dc
1cc304c3
1d935664
98ac388c
516c0c33
71ec082b
05946087
ffc4325c
02d3540c
f04ed23c
a3c3740c
74dcdae4
a830000d
a3c3742c
14dcdae4
a850000d
a3c3744c
b4dcdae4
686c000c
a2c3546c
54dc3ae4
4e57000c
03e432c3
000c04dc
606c09c3
111c2006
31830004
32dc6007
5b3c000b
05c30e00
f6bc3fe6
788c09e2
185163f2
78ac0473
0a9443e4
78af702c
10c318cc
179441e4
58cf4006
4c2c0293
42e40213
102c0c94
38cc0c2f
42e421c3
78cf0294
000678cc
00b30c2f
482c32c3
009351f2
7fe5788c
05c3788f
09e476bc
20071053
29c39f94
0006686c
0004011c
60073083
3c2f7894
64d278ac
ec2f78cc
f8af0053
788cf8cf
788f6025
106c401c
0000411c
6cac700c
6c546007
16c308c3
30c33664
60073264
700c6554
68d26cec
17c308c3
366426c3
326430c3
f8ac64f2
38af3c2c
7fe5788c
301c788f
311c106c
6c0c0000
46f24c89
d8ec08d3
94dc62e4
7decffbf
540c6ef7
03946087
01134f37
142c4f37
344c0f77
546c2fb7
39c34ff7
31c32c6c
011c0006
30830004
2b946007
09c37ccc
4c00002c
e08c313c
49a06212
4c2f39c3
000631c3
0002011c
65d23083
0010323c
642f19c3
10002f3c
f64e323c
07946087
9f5c4037
0bc30027
00f32006
40377f0c
00279f5c
13c30bc3
6e572cc3
0a0b3abc
66bc07c3
00930a40
3fe5902c
4096ef33
0f56fc76
00000804
0136f016
50c3f496
005c71c3
10c304c1
04c9055c
40ac303c
04d1155c
81ac313c
04d9255c
c1ac823c
10c31689
303c16a9
36c940ac
81ac313c
423c56e9
38c3c1ac
06e4035c
02c01f3c
0b948087
60064706
0a4e5abc
54dc0007
62d7002a
11f38def
60064706
0a4e5abc
b4dc0007
62d70029
0def00c6
370942d7
372901c3
402c313c
303c1749
376981ac
c1ac313c
42d76a0f
10c31789
303c17a9
37c940ac
81ac313c
303c17e9
6a2fc1ac
155c42d7
01c30101
0109155c
402c313c
0111055c
81ac303c
0119155c
c1ac313c
42d76a4f
0121055c
055c10c3
303c0129
155c40ac
313c0131
055c81ac
303c0139
6a6fc1ac
155c42d7
01c30a21
0a29155c
402c313c
0a31055c
81ac303c
0a39155c
c1ac313c
0a8f0c4c
155c42d7
01c30a21
0a29155c
402c313c
0a31055c
81ac303c
0a39155c
c1ac313c
0aaf0c6c
155c42d7
01c30a21
0a29155c
402c313c
0a31055c
81ac303c
0a39155c
c1ac313c
0acf0c8c
155c42d7
01c30a21
0a29155c
402c313c
0a31055c
81ac303c
0a39155c
c1ac313c
0aef0cac
155c42d7
01c30181
0189155c
402c313c
0191055c
81ac303c
0199155c
c1ac313c
42d768ef
01a1055c
055c10c3
303c01a9
155c40ac
313c01b1
055c81ac
303c01b9
690fc1ac
696c42d7
698f6385
238662d7
62d72ccf
7589cd6c
75a903c3
402c233c
0141055c
055c10c3
303c0149
155c40ac
313c0151
055c81ac
303c0159
323cc1ac
780f81ac
155cf82f
21c30201
0209155c
412c313c
0211255c
81ac323c
0219055c
c1ac303c
17946067
584f4006
03c1055c
055c10c3
303c03c9
155c40ac
313c03d1
255c81ac
323c03d9
0006c1ac
7002011c
049330a3
0241155c
155c21c3
313c0249
255c412c
323c0251
055c81ac
303c0259
784fc1ac
03c1155c
155c21c3
313c03c9
255c412c
323c03d1
055c81ac
303c03d9
2006c1ac
7012111c
786f31a3
02c35689
323c56a9
16c9402c
81ac303c
313c36e9
42d7c1ac
15946087
6d2c68ec
fd80233c
3f5c42b7
760d0141
ffff241c
483242b7
1f5c4277
362d0121
564d4006
0293566d
6d2c68ec
fc40133c
2f5c2237
560d0101
ffff141c
28322237
0f5c21f7
162d00e1
364d2006
255c366d
02c303c1
03c9255c
402c323c
03d1055c
81ac303c
03d9155c
c1ac213c
560941b7
562902c3
402c323c
303c1649
366981ac
c1ac313c
02c34197
183530e4
00c11f5c
4197360d
420b323c
3f5c6177
762d00a1
103c0197
2137440b
00811f5c
4197364d
40f75832
00613f5c
0006766d
3609188f
362921c3
412c313c
323c5649
166981ac
c1ac103c
211c4006
12a30204
323c580c
3203818c
418c223c
ffff001c
ff00011c
68323083
780f3203
323c582c
3203818c
418c223c
68323083
782f3203
323c584c
3203818c
418c223c
68323083
784f3203
323c586c
3203818c
418c223c
68323083
786f3203
818c313c
213c3103
3083418c
32036832
101c78af
111c0101
38cf0001
02c35689
323c56a9
16c9402c
81ac303c
313c36e9
6087c1ac
055c1394
10c30181
0189055c
40ac303c
0191155c
81ac313c
0199255c
c1ac323c
0140733c
055c0253
10c30a21
0a29055c
40ac303c
0a31155c
81ac313c
0a39255c
c1ac323c
0080733c
88cc42d7
0180353c
02c36037
24c320c6
38bc37c3
30e30a3f
800c233c
818c323c
223c3203
001c418c
011cffff
3083ff00
32036832
3689788f
36a921c3
412c313c
323c56c9
16e981ac
c1ac303c
608742d7
055c5594
10c30181
0189055c
40ac303c
0191155c
81ac313c
0199055c
c1ac303c
370968ef
372921c3
412c313c
323c5749
176981ac
c1ac203c
04e1155c
155c01c3
313c04e9
055c402c
303c04f1
155c81ac
413c04f9
055cc1ac
10c30501
0509055c
40ac303c
0511155c
81ac313c
0519055c
c1ac303c
20066037
0006111c
055c2077
10c30521
0529055c
40ac303c
0531155c
81ac313c
0539055c
c1ac303c
08c360b7
34c322d7
0a22a0bc
155c0453
01c30a21
0a29155c
402c313c
0a31055c
81ac303c
0a39155c
c1ac313c
42d76b0f
106c301c
0000311c
a8cc6c0c
005c08c3
003731a4
08c38e4c
40c612c3
466435c3
80760c96
08040f56
0336f016
40c3f796
0f3c71c3
256c0100
b0bc4286
045c08cb
10c30201
0209045c
40ac303c
0211145c
81ac313c
0219245c
c1ac523c
09b4a067
c00661d7
0004611c
60073683
000b72dc
00e48f5c
383c2157
233ce08c
7ccc100c
60f76d20
0241045c
045c20c3
303c0249
245c412c
323c0251
645c81ac
263c0259
045cc1ac
60c303a1
03a9045c
432c303c
03b1645c
81ac363c
03b9045c
c1ac603c
600760d7
0f5c1f94
30c30061
6026c2f2
60b73264
12e463d2
00973a54
35940007
60076520
3f5c3274
03c30041
6ca07900
02f46007
203c0026
40770016
00212f5c
c0070473
65202254
0a746007
60a01900
06f46007
93c360d7
09e49184
313c1834
6d20fff0
6c0000d7
0f746007
79000006
20d76ca0
60076ca0
00260274
0016603c
2f5cc037
00930001
00534026
38c34006
011c0006
30830004
28546007
0994a067
c00638c3
0010611c
60073683
000dd2dc
a06744d2
000d94dc
0221045c
045c10c3
303c0229
145c40ac
313c0231
645c81ac
263c0239
6197c1ac
045432e4
42dca067
04c3000c
0a1316bc
400717f3
07c31754
0a4066bc
0221145c
145c21c3
313c0229
245c412c
323c0231
04c381ac
0239645c
c1ac163c
0a0cd6bc
a0c71553
a0c74b54
a08709b4
a0871654
a0671fb4
000824dc
a1070153
a1076754
a1275314
a1677554
09137894
1f3c04c3
22bc0100
00d30a18
1f3c04c3
76bc0100
04c30a16
00bc17c3
50c30a37
6f3c0cf3
04c30100
b4bc16c3
50c30a47
106c801c
0000811c
28c307f2
6c4c680c
13946007
04c30a93
00bc17c3
50c30a37
16c304c3
0a14fcbc
4ebc04c3
68c30a1a
6c4c780c
44546007
366404c3
04c30833
01001f3c
0a47b4bc
39540007
17c304c3
0a3700bc
04c350c3
0a1a4ebc
04c30633
01001f3c
0a15c6bc
6f3c0553
04c30100
b4bc16c3
00070a47
04c32254
00bc17c3
50c30a37
16c304c3
0a54c0bc
6f3c0333
04c30100
b4bc16c3
00070a47
04c31054
00bc17c3
50c30a37
16c304c3
0a561abc
04c300f3
01001f3c
0a145cbc
61d7a006
011c0006
30830020
13546007
08a1145c
145c21c3
313c08a9
245c412c
323c08b1
645c81ac
363c08b9
63d2c1ac
366404c3
07c3a4f2
0a4066bc
c0760996
08040f56
3f36f016
50c3ca96
d2c361c3
10c30289
303c16a9
36c940ac
81ac313c
123c56e9
2087c1ac
455c1394
04c30181
0189455c
402c343c
0191055c
81ac303c
0199255c
c1ac323c
0140c33c
20c70333
005634dc
0a21455c
455c04c3
343c0a29
055c402c
303c0a31
455c81ac
243c0a39
6849c1ac
04dc6087
c23c0055
b53c0080
39ef0180
0246784c
aaaa101c
aaaa111c
32e421c3
005424dc
f5244e24
0701455c
455c04c3
343c0709
055c402c
303c0711
155c81ac
313c0719
6bf2c1ac
4004323c
60070486
0052a2dc
0486f324
0005269c
0201455c
455c04c3
343c0209
055c402c
303c0211
155c81ac
313c0219
7f65c1ac
0400241c
07356027
40070706
0050e2dc
2bd3f324
04c1055c
055c10c3
303c04c9
155c40ac
313c04d1
455c81ac
a43c04d9
42d2c1ac
055cf324
10c30181
0189055c
40ac303c
0191155c
81ac313c
0199255c
c1ac323c
455c78ef
04c301a1
01a9455c
402c343c
01b1055c
81ac303c
01b9155c
c1ac313c
796c790f
fec0433c
78cc996f
78cf6285
03c37589
233c75a9
055c402c
10c30141
0149055c
40ac303c
0151155c
81ac313c
0159055c
c1ac303c
81ac323c
155c700f
21c30241
0249155c
412c313c
0251255c
81ac323c
0259055c
c1ac303c
155c704f
21c303c1
03c9155c
412c313c
03d1255c
81ac323c
03d9055c
c1ac303c
111c2006
31a35018
4006706f
055c508f
10c30241
0249055c
40ac303c
0251155c
81ac313c
0259255c
c1ac023c
3f5c0d77
355c06a1
103c0265
2d37420b
06812f5c
026d255c
033c6d57
0cf7440b
06610f5c
0275055c
38322d57
2f5c2cb7
255c0641
055c027d
10c303c1
03c9055c
40ac303c
03d1155c
81ac313c
03d9255c
c1ac023c
3f5c0c77
355c0621
103c03e5
2c37420b
06012f5c
03ed255c
033c6c57
0bf7440b
05e10f5c
03f5055c
38322c57
2f5c2bb7
255c05c1
301c03fd
311c1108
0c090000
0285055c
155c2c29
4c49028d
0295255c
055c0c69
500c029d
818c323c
223c3203
101c418c
111cffff
3183ff00
32036832
504c700f
818c323c
223c3203
3183418c
32036832
506c704f
818c323c
223c3203
3183418c
32036832
508c706f
818c323c
223c3203
3183418c
32036832
8a3c708f
155c0e00
21c30221
0229155c
412c313c
0231255c
81ac323c
0239055c
c1ac703c
818c373c
273c3703
101c418c
111cffff
3183ff00
32036832
78cc702f
0007bf5c
20c606c3
3cc323c3
0a3f38bc
93c330e3
08c39364
f6bc3fe6
055c09e2
10c30221
0229055c
40ac303c
0231155c
81ac313c
0239255c
c1ac323c
055473e4
76bc08c3
f81309e4
0201155c
155c21c3
313c0209
255c412c
323c0211
055c81ac
303c0219
7f65c1ac
06356027
76bc08c3
070609e4
4e247593
18ccf524
033c7c00
0b77fec0
05a11f5c
0225155c
420b003c
1f5c0b37
155c0581
6b57022d
440b033c
0f5c0af7
055c0561
2b570235
2ab73832
05413f5c
023d355c
4004323c
f32462d2
800c293c
818c323c
223c3203
001c418c
011cffff
3083ff00
32036832
155c708f
21c305c1
05c9155c
412c313c
05d1255c
81ac323c
05d9455c
c1ac243c
05a1055c
055c10c3
303c05a9
155c40ac
313c05b1
455c81ac
343c05b9
23e4c1ac
002581dc
05e1155c
155c21c3
313c05e9
255c412c
323c05f1
455c81ac
043c05f9
0a77c1ac
0ff4163c
363c21b7
6177408c
808c063c
263c0137
40f7c08c
60076a57
455c2254
04c30601
0609455c
402c343c
0611055c
81ac303c
0619155c
c1ac313c
2f5ccc4f
255c00c1
3f5c0605
355c00a1
4f5c060d
455c0081
0f5c0615
055c0061
0ed3061d
00c11f5c
05e5155c
32c34157
00ff341c
4f5c6a37
455c0501
011705ed
141c10c3
29f700ff
04e12f5c
05f5255c
00613f5c
05fd355c
00c14f5c
0605455c
05010f5c
060d055c
04e11f5c
0615155c
00612f5c
061d255c
0641455c
455c04c3
343c0649
055c402c
303c0651
155c81ac
213c0659
49b7c1ac
04c12f5c
0625255c
433c6997
8977420b
04a14f5c
062d455c
103c0997
2937440b
04811f5c
0635155c
58324997
3f5c48f7
355c0461
4f5c063d
455c0521
0f5c0665
055c0521
1f5c066d
155c0521
2f5c0675
255c0521
3f5c067d
355c0521
4f5c0325
455c0521
0f5c032d
055c0521
1f5c0335
155c0521
201c033d
211ceeee
584feeee
05c1455c
455c04c3
343c05c9
055c402c
303c05d1
155c81ac
313c05d9
433cc1ac
88b70010
04410f5c
05c5055c
420b243c
3f5c4877
355c0421
043c05cd
0837440b
04011f5c
05d5155c
58324897
3f5c47f7
355c03e1
455c05dd
04c30321
0329455c
402c343c
0331055c
81ac303c
0339155c
c1ac313c
6d0058cc
fec0033c
1f5c07b7
155c03c1
303c0325
6777420b
03a14f5c
032d455c
440b103c
2f5c2737
255c0381
67970335
66f77832
03614f5c
033d455c
0401055c
055c10c3
303c0409
155c40ac
313c0411
255c81ac
323c0419
033cc1ac
06b70010
03411f5c
0405155c
420b303c
4f5c6677
455c0321
103c040d
2637440b
03012f5c
0415255c
78326697
4f5c65f7
455c02e1
055c041d
10c30421
0429055c
40ac303c
0431155c
81ac313c
0439255c
c1ac323c
6e0098cc
fec0133c
2f5c25b7
255c02c1
413c0425
8577420b
02a10f5c
042d055c
440b213c
3f5c4537
355c0281
85970435
84f79832
02610f5c
043d055c
21c33689
313c36a9
56c9412c
81ac323c
343c96e9
3709c1ac
17495729
6087f769
323c4094
203c40ac
055c81ac
10c304e1
04e9055c
40ac303c
04f1155c
81ac313c
04f9055c
c1ac403c
0501155c
155c01c3
313c0509
055c402c
303c0511
155c81ac
313c0519
6037c1ac
311c6006
60770006
0521055c
055c10c3
303c0529
155c40ac
313c0531
055c81ac
303c0539
60b7c1ac
16c30ac3
c12c273c
a0bc34c3
13130a22
40ac323c
81ac303c
c1ac373c
37897a0f
37a921c3
412c313c
323c57c9
97e981ac
c1ac343c
055c7a2f
10c30101
0109055c
40ac303c
0111155c
81ac313c
0119255c
c1ac323c
455c7a4f
04c30121
0129455c
402c343c
0131055c
81ac303c
0139155c
c1ac313c
255c7a6f
42c30a21
0a29255c
422c323c
0a31455c
81ac343c
0a39055c
c1ac303c
3a8f2c4c
0a21255c
255c42c3
323c0a29
455c422c
343c0a31
055c81ac
303c0a39
2c6cc1ac
255c3aaf
42c30a21
0a29255c
422c323c
0a31455c
81ac343c
0a39055c
c1ac303c
3acf2c8c
0a21255c
255c42c3
323c0a29
455c422c
343c0a31
055c81ac
303c0a39
2cacc1ac
255c3aef
42c30a21
0a29255c
422c323c
0a31455c
81ac343c
0a39055c
c1ac303c
301c7b0f
311c106c
6c0c0000
1ac3b8cc
31a4115c
8e4c2037
16c30ac3
35c340c6
08c34664
09e476bc
20330006
40072dc3
000a02dc
11b4401c
0000411c
3a3c500c
23e414c0
000962dc
07c1155c
155c01c3
313c07c9
055c402c
303c07d1
155c81ac
313c07d9
6007c1ac
255c3954
42c30221
0229255c
422c323c
0231455c
81ac343c
0239055c
c1ac303c
38cc6285
64b76ca0
02412f5c
0225255c
420b433c
0f5c8477
055c0221
2497022d
440b213c
2f5c4437
255c0201
64970235
63f77832
01e14f5c
023d455c
7d8578cc
796c78cf
796f6285
76bc08c3
080609e4
cbef1553
07c1055c
055c10c3
303c07c9
155c40ac
313c07d1
255c81ac
323c07d9
133cc1ac
23b70010
01c12f5c
07c5255c
420b013c
1f5c0377
155c01a1
439707cd
440b323c
3f5c6337
355c0181
039707d5
02f71832
01611f5c
07dd155c
0007df5c
0f40053c
209c101c
0014111c
38c325c3
0a5776bc
335c700c
67d20424
7d8578cc
796c78cf
796f6285
11b4301c
0000311c
035c6c0c
0bf30424
0221255c
255c42c3
323c0229
455c422c
343c0231
055c81ac
303c0239
6285c1ac
6ca038cc
2f5c62b7
255c0141
433c0225
8277420b
01210f5c
022d055c
213c2297
4237440b
01012f5c
0235255c
78326297
4f5c61f7
455c00e1
78cc023d
78cf7d85
6285796c
055c796f
10c305c1
05c9055c
40ac303c
05d1155c
81ac313c
05d9455c
c1ac243c
05a1055c
055c10c3
303c05a9
155c40ac
313c05b1
455c81ac
343c05b9
23e4c1ac
08c30634
09e476bc
00f30726
76bc08c3
092609e4
0a060053
fc763696
08040f56
40c37016
40cc51c3
13e432c3
20073134
205c2f54
6100fd53
fd6e135c
6ca060cc
616c60cf
616f6285
618c216c
56e4cca0
04e41535
318f0394
406c0193
6006506f
201c606f
211caaaa
404faaaa
0a4066bc
106cb720
e994a007
04e40113
6ea00494
0073718f
616f6680
7d85716c
0e56716f
00000804
40c37016
13e460cc
aca02734
301ca0cf
311c106c
6c0c0000
62d26d0c
04c33664
818c0333
7120416c
35e4206c
6a200415
01f3b580
618f6a80
606f6006
501c2ad2
511caaaa
a44faaaa
66bc01c3
00930a40
000701c3
0e56e794
00000804
3f36f016
50c38f96
056c3af7
206c1bb7
313c0030
233ce08c
9ad7100c
b3c370cc
0bc3b2a4
1bf70884
400631c3
0001211c
60073283
3f5c2454
355c0de1
603c02a5
dab7420b
0d417f5c
02ad755c
440b103c
2f5c3a77
255c0d21
7bd702b5
7a377832
0d014f5c
02bd455c
655cc026
e00602c5
02cd755c
02d5755c
02dd755c
00070bc3
155c5294
21c30201
0209155c
412c313c
0211255c
81ac323c
0219455c
c1ac343c
04dc60a7
755c007e
07c30541
0549755c
402c373c
0551055c
81ac303c
0559155c
c1ac313c
e4dc6007
255c007c
42c30241
0249255c
422c323c
0251455c
81ac343c
0259655c
c1ac363c
5c2cfb97
a2dc32e4
7fe5007b
62dc32e4
255c007b
42c30221
0229255c
422c323c
0231455c
81ac343c
655c05c3
163c0239
d6bcc1ac
0bc30a0c
0007a49c
fad70006
155c1c2f
21c30581
0589155c
412c313c
0591255c
81ac323c
0599455c
c1ac043c
416c0ad2
c82c60cc
686c2f00
62127c32
021325a0
0241755c
755c17c3
373c0249
155c40ac
313c0251
255c81ac
123c0259
7b97c1ac
455c4c2c
64c30241
0249455c
432c343c
0251655c
81ac363c
0259755c
c1ac473c
84dc24e4
12e4000c
000c54dc
bbbb101c
bbbb111c
3c2ffad7
00ff741c
7ad7e137
60f76832
90329ad7
dad780b7
c077d832
14540007
e04ffad7
00810f5c
0585055c
00611f5c
058d155c
00412f5c
0595255c
00213f5c
059d355c
4f5c0713
455c0081
c0d70565
741c76c3
f9f700ff
0ce10f5c
056d055c
21c32097
00ff241c
3f5c59b7
355c0cc1
4f5c0575
455c0021
6f5c057d
655c0081
70c30585
058d755c
055c03c3
14c30595
059d155c
1108301c
0000311c
255c4c09
8c290285
028d455c
655ccc49
ec690295
029d755c
0541055c
055c10c3
303c0549
155c40ac
313c0551
255c81ac
323c0559
633cc1ac
d9770010
0ca17f5c
0545755c
420b163c
2f5c3937
255c0c81
463c054d
98f7440b
0c616f5c
0555655c
f832f957
0f5cf8b7
055c0c41
201c055d
211ceeee
3ad7eeee
7b97444f
78776c6c
0c214f5c
02e5455c
ffff341c
68327877
7f5c7837
755c0c01
000602ed
02f5055c
02fd055c
0de11f5c
0245155c
323c5bd7
77f7420b
0be13f5c
024d355c
643c9bd7
d7b7440b
0bc16f5c
0255655c
f832fbd7
0f5cf777
055c0ba1
901c025d
c9c30001
155c6d73
21c30561
0569155c
412c313c
0571255c
81ac323c
0579755c
c1ac673c
34dcc007
84e4000a
48a42b15
14c31ad7
0a3698bc
1f5cb4a4
155c0de1
5bd70245
420b323c
3f5c7737
355c0b81
9bd7024d
440b643c
6f5cd6f7
655c0b61
fbd70255
f6b7f832
0b410f5c
025d055c
bbbb201c
bbbb211c
442f3ad7
0001901c
455c0293
74c30221
0229455c
43ac343c
0231755c
81ac373c
255c05c3
123c0239
d6bcc1ac
96c30a0c
7ad7c9c3
441c43c3
967700ff
0b216f5c
0565655c
073cfad7
1637420b
0b010f5c
056d055c
213c3ad7
55f7440b
0ae12f5c
0575255c
78327ad7
4f5c75b7
455c0ac1
655c057d
70c30585
058d755c
055c02c3
14c30595
059d155c
255c4026
60060545
054d355c
0555355c
055d355c
1108301c
0000311c
455c8c09
cc290285
028d655c
755cec49
0c690295
029d055c
eeee201c
eeee211c
444f3ad7
6c6c7b97
4f5c7577
455c0aa1
341c02e5
7577ffff
75376832
0a817f5c
02ed755c
055c0006
055c02f5
571302fd
2c1584e4
1ad748a4
98bc14c3
b4a40a36
2f5c8484
255c0de1
7bd70245
420b433c
4f5c94f7
455c0a61
dbd7024d
440b763c
7f5cf4b7
755c0a41
1bd70255
14771832
0a211f5c
025d155c
bbbb301c
bbbb311c
682f5ad7
0001901c
901c0353
c9c30000
16f484e4
0221755c
755c07c3
373c0229
055c402c
303c0231
05c381ac
0239255c
c1ac123c
0a0cd6bc
0000901c
455cc9c3
64c30561
0569455c
432c343c
0571655c
81ac363c
0579755c
c1ac673c
0000a01c
001c3073
011ceeee
10c3eeee
039461e4
2fb3c006
ec2c796c
5e0098cc
7c326c6c
49a06212
d2a4d8c3
0000d31c
0016b8dc
9da07bd7
b8dc8007
38c30016
20072fa0
1bd72d74
60076820
155c2974
21c30241
0249155c
412c313c
0251255c
81ac323c
0259455c
c1ac343c
79a068c3
87dc6007
055c0055
10c30221
0229055c
40ac303c
0231155c
81ac313c
255c05c3
123c0239
d6bcc1ac
449c0a0c
08c30005
60077c20
000cf3dc
61201bd7
f3dc6007
984c000b
aaaa101c
aaaa111c
055c384f
10c30541
0549055c
40ac303c
0551155c
81ac313c
0559055c
c1ac303c
fff0033c
1f5c1437
155c0a01
003c0545
13f7420b
09e11f5c
054d155c
033c7417
13b7440b
09c10f5c
0555055c
38323417
3f5c3377
355c09a1
06c3055d
66bc4037
655c0a40
06c30441
0449655c
402c363c
0451055c
81ac303c
0459155c
c1ac313c
fff0033c
1f5c1337
155c0981
603c0445
d2f7420b
09610f5c
044d055c
313c3317
72b7440b
09413f5c
0455355c
d832d317
0f5cd277
055c0921
155c045d
61c30461
0469155c
432c313c
0471655c
81ac363c
0479055c
c1ac303c
40176f80
72376d20
09011f5c
0465155c
420b633c
0f5cd1f7
055c08e1
3217046d
440b313c
3f5c71b7
355c08c1
d2170475
d177d832
08a10f5c
047d055c
03c1155c
155c61c3
313c03c9
655c432c
363c03d1
055c81ac
303c03d9
6fa0c1ac
71376d00
08811f5c
03c5155c
420b333c
6f5c70f7
655c0861
f11703cd
440b073c
0f5c10b7
055c0841
311703d5
30773832
08212f5c
03dd255c
0e1364c3
68201bd7
08f46007
5bd71ad7
d2bc2ba0
b4840a36
20070d13
9bd76374
600773a0
08c35ff4
06c38820
d2bc14c3
155c0a36
21c30461
0469155c
412c313c
0471255c
81ac323c
0479755c
c1ac373c
df5cd384
1f5c0807
155c0801
3d3c0465
6ff7420b
07e13f5c
046d355c
440b0d3c
0f5c0fb7
055c07c1
1dc30475
2f773832
07a12f5c
047d255c
03c1755c
755c07c3
373c03c9
055c402c
303c03d1
155c81ac
313c03d9
7180c1ac
2f5c6f37
255c0781
433c03c5
8ef7420b
07617f5c
03cd755c
103c0f17
2eb7440b
07411f5c
03d5155c
58324f17
3f5c4e77
355c0721
a6c303dd
c007d84c
ffe7d4dc
80074ac3
7f5c1d94
755c0d61
1ad70565
420b103c
1f5c2e37
155c0701
5ad7056d
440b323c
3f5c6df7
355c06e1
9ad70575
8db79832
06c17f5c
057d755c
3ad70093
204f0ac3
2394c007
0d612f5c
0585255c
433c7ad7
8d77420b
06a14f5c
058d455c
763cdad7
ed37440b
06817f5c
0595755c
18321ad7
1f5c0cf7
155c0661
301c059d
311ceeee
5ad7eeee
0073684f
d04f9ad7
0541655c
655c76c3
363c0549
755c43ac
373c0551
055c81ac
303c0559
233cc1ac
4cb70010
06413f5c
0545355c
420b623c
7f5ccc77
755c0621
123c054d
2c37440b
06012f5c
0555255c
78326c97
4f5c6bf7
455c05e1
655c055d
76c30561
0569655c
43ac363c
0571755c
81ac373c
0579055c
c1ac103c
0241255c
255c42c3
323c0249
455c422c
343c0251
655c81ac
463c0259
656cc1ac
0c2ccc6c
702044cc
30746007
363c4800
6212e08c
7c3769a0
60076e20
2f5c2ff4
255c0e01
7c170245
420b433c
4f5c8bb7
455c05c1
dc17024d
440b763c
7f5ceb77
755c05a1
1c170255
0b371832
05812f5c
025d255c
0001c21c
bbbb301c
bbbb311c
9c17642f
0001901c
642c0133
bbbb601c
bbbb611c
37e476c3
244c0b94
eeee001c
eeee011c
12e420c3
20070354
455cb994
64c30441
0449455c
432c343c
0451655c
81ac363c
0459755c
c1ac373c
0010133c
2f5c2af7
255c0561
413c0445
8ab7420b
05416f5c
044d655c
440b013c
1f5c0a77
155c0521
4ad70455
4a375832
05013f5c
045d355c
0461455c
455c64c3
343c0469
655c432c
363c0471
755c81ac
373c0479
0bc3c1ac
09f70180
04e11f5c
0465155c
420b303c
4f5c69b7
455c04c1
703c046d
e977440b
04a10f5c
0475055c
383229d7
2f5c2937
255c0481
455c047d
64c303c1
03c9455c
432c343c
03d1655c
81ac363c
03d9755c
c1ac373c
4c34b3e4
13c33ba4
2f5c7b37
255c0d81
433c03c5
88f7420b
04616f5c
03cd655c
440b013c
0f5c08b7
055c0441
383203d5
2f5c2877
255c0421
455c03dd
64c303a1
03a9455c
432c343c
03b1655c
81ac363c
03b9755c
c1ac073c
083770c3
20c31b17
27e417c3
3f5c2435
355c0401
673c03c5
c7f7420b
03e17f5c
03cd755c
440b113c
2f5c27b7
255c03c1
681703d5
67777832
03a14f5c
03dd455c
c0060153
03c5655c
03cd655c
03d5655c
03dd655c
03e1755c
755c07c3
373c03e9
055c402c
303c03f1
155c81ac
313c03f9
b3e4c1ac
3ba41d34
6f5c6737
655c0381
033c03e5
06f7420b
03611f5c
03ed155c
440b333c
4f5c66b7
455c0341
c71703f5
c677d832
03217f5c
03fd755c
00060153
03e5055c
03ed055c
03f5055c
03fd055c
0ec0453c
155c3173
21c30561
0569155c
412c313c
0571255c
81ac323c
0579655c
c1ac163c
0541755c
755c07c3
373c0549
055c402c
303c0551
255c81ac
323c0559
6027c1ac
e0061394
0565755c
056d755c
0575755c
057d755c
0585755c
058d755c
0595755c
059d755c
050901b3
0565055c
255c4529
6549056d
0575355c
655cc569
701c057d
711caaaa
e44faaaa
042f0006
0541255c
255c62c3
323c0549
655c432c
363c0551
755c81ac
373c0559
233cc1ac
4637fff0
03013f5c
0545355c
420b723c
0f5ce5f7
055c02e1
323c054d
65b7440b
02c16f5c
0555655c
f832e617
0f5ce577
055c02a1
456c055d
686c5bb7
233c7c32
db97100c
656f7900
6d2064cc
755c64cf
07c30761
0769755c
402c373c
0771055c
81ac303c
0779255c
c1ac323c
2c0f6fec
03c1655c
655c76c3
363c03c9
755c43ac
373c03d1
055c81ac
303c03d9
44ccc1ac
7b776d00
0da13f5c
03c5355c
763cdb57
e537420b
02817f5c
03cd755c
103c1b57
24f7440b
02611f5c
03d5155c
58325b57
3f5c44b7
355c0241
655c03dd
76c303a1
03a9655c
43ac363c
03b1755c
81ac373c
03b9055c
c1ac103c
247701c3
31c33b57
30e420c3
6f5c1a35
655c0221
003c03c5
0437420b
02011f5c
03cd155c
440b323c
3f5c63f7
355c01e1
c45703d5
c3b7d832
01c17f5c
03dd755c
0781055c
055c10c3
303c0789
155c40ac
313c0791
255c81ac
323c0799
733cc1ac
e377fff0
01a10f5c
0785055c
420b273c
3f5c4337
355c0181
773c078d
e2f7440b
01610f5c
0795055c
38322357
2f5c22b7
255c0141
655c079d
76c303c1
03c9655c
43ac363c
03d1755c
81ac373c
03d9055c
c1ac203c
03e1155c
155c61c3
313c03e9
655c432c
363c03f1
755c81ac
373c03f9
49a0c1ac
03a1055c
055c10c3
303c03a9
155c40ac
313c03b1
655c81ac
363c03b9
6132c1ac
401423e4
0541055c
055c10c3
303c0549
155c40ac
313c0551
255c81ac
323c0559
6007c1ac
db972f94
e006786c
0001711c
60073783
055c2794
10c30201
0209055c
40ac303c
0211155c
81ac313c
0219255c
c1ac323c
169460a7
e00779c3
055c1354
10c30221
0229055c
40ac303c
0231155c
81ac313c
255c05c3
123c0239
d6bcc1ac
c21c0a0c
04c3ffff
38bc2006
3cc30a57
13546007
0761655c
655c76c3
363c0769
755c43ac
373c0771
055c81ac
303c0779
6007c1ac
ffe634dc
200719c3
0009d2dc
0961255c
255c42c3
323c0969
455c422c
343c0971
655c81ac
363c0979
6007c1ac
02f31594
ffffc21c
0961755c
755c07c3
373c0969
055c402c
303c0971
155c81ac
313c0979
05c3c1ac
2cc33664
eb944007
106c301c
0000311c
6c0c6c0c
40074da9
455c6b54
64c30201
0209455c
432c343c
0211655c
81ac363c
0219755c
c1ac373c
5a9460a7
246c3b97
311c6006
13830001
20072277
455c5194
64c30341
0349455c
432c343c
0351655c
81ac363c
0359755c
c1ac373c
211432e4
155c2026
2f5c0345
255c0121
32c3034d
0355355c
455c42c3
655c035d
76c30221
0229655c
43ac363c
0231755c
81ac373c
255c05c3
123c0239
d6bcc1ac
04130a0c
0010633c
7f5cc237
755c0101
163c0345
21f7420b
00e12f5c
034d255c
440b463c
6f5c81b7
655c00c1
e2170355
e177f832
00a10f5c
035d055c
00060073
00260053
fc767196
08040f56
1f36f016
a0c3ff96
52c361c3
e2d703c3
0116313c
0b0d333c
b33c7fe5
1bc3f88c
c74726f2
4bc30454
2d94c0c7
e3f202d2
22330026
7a00800b
6c80202b
6d005c0b
2e009c2b
69ec2ac3
0c9460c7
373c4046
83c3259d
259d303c
18848384
41074025
6680f794
808c233c
ffff341c
233c6d00
341c808c
4d00ffff
408c323c
41ac423c
ffff441c
400c0ac3
0046363c
0b0d333c
7f3233c4
84dc4027
60070008
000852dc
f6809a3c
325c29c3
801c0404
001c0000
011ccccc
10c30000
2a9431e4
0424325c
808c233c
ffff341c
3ac34d00
0106ed6c
25f21bc3
c0c70bc3
02860294
808c323c
ffff241c
13e36980
ffff141c
088c303c
00b34006
259d673c
40252700
fb1423e4
5d806112
0ac39080
b42000cc
183c1113
213c0010
313c0014
333c088c
6d000067
29c360c5
359d223c
400646f2
b93c02c3
00b32000
20a781c3
ff13eb94
088c703c
0014603c
0067373c
133c6f00
39c30060
159d133c
63542007
6ac30bf2
1bc3596c
53e46520
353c1b34
2980fff0
373c02f3
6f000037
69c36085
3a1d263c
0001831c
313c0594
2980fff0
28800053
ffff821c
323c00b3
9180013f
21e4bfc5
0025fb14
cd9400c7
40070793
60072e94
3a3c2c54
035cfa80
ba3c0293
73c31a80
62c380c3
03d39bc3
1ac3cbf2
19c3456c
1bc36520
103453e4
fff0353c
5c4c00f3
831c7ccb
02940001
29807fe5
323c00b3
9180013f
21e4bfc5
821cfb14
c025ffff
60e4e105
01b3e214
416c0ac3
fff0353c
00b32980
013f323c
bfc59180
fb1421e4
0b94a027
00403f3c
033c080b
2006ff6e
2f5c2c2d
91000013
808c343c
ffff441c
233c7180
341c808c
4d00ffff
408c323c
41ac323c
036403c3
f8760196
08040f56
40c3f016
106c301c
0000311c
6c8c6c0c
62546007
30c33664
60273264
0cb35d94
300c704c
aaaa201c
aaaa211c
30e402c3
20070f54
640c5c54
434b201c
5041211c
30e402c3
64cc5494
64cf6025
d06c0a13
056cf524
34540007
03e4638c
60060494
00f3656f
438c656f
6baf63ac
4f8f63ac
7fe5658c
4006658f
7c0c434f
7c0f6025
f324a2d2
706f6006
708f702f
712c70cf
6d0043cc
718f716f
70ef6006
201c710f
211caaaa
504faaaa
01c5345c
51ef4006
8c0f63ec
0427205c
09f102bc
7fe60173
04ec704f
84ef106f
6025644c
a2d2644f
46c3f324
6e240113
4004533c
1250701c
0000711c
9d948007
00530006
0f5600e6
00000804
106c301c
0000311c
6d6c6c0c
366401c3
00000804
0136f016
41c370c3
79a9c56c
798983c3
442c533c
0787323c
1070801c
0000811c
480c28c3
4c4c6d00
531c44ef
08540800
86dd201c
0000211c
53e432c3
716c0c94
716f61c5
7e4570cc
07c370cf
3abc14c3
04130a07
0806531c
363c0a94
656f00e0
7e4564cc
28bc64cf
02930a05
8035201c
0000211c
53e432c3
363c0a94
656f00e0
7e4564cc
0cbc64cf
00930a57
66bc01c3
80760a40
08040f56
0736f016
2006fe96
20d02077
a0ec202f
800cd4e9
3d548267
1070301c
0000311c
640c2c0c
646c69d2
069439e4
a01c644c
35e40000
21c30e54
3c4e323c
60546007
39e4686c
684c5d94
5a9435e4
0001a01c
0db480e7
78348087
54548027
74548007
6c548047
b4dc8067
0d730012
12dc8147
81470012
810708b4
000d02dc
f4dc8127
1df30011
d2dc8247
82670011
001184dc
1070301c
0000311c
680c4c0c
65d213c3
60076bcc
20262d94
0787513c
6ae16026
1070601c
0000611c
6e80780c
780c2c2f
80ec6e80
780c8c4f
2c716e80
10e8401c
0000411c
7f5cf009
10290035
003d0f5c
ee80780c
00400f3c
09f7eabc
780c1c8f
043cae80
eabc0020
14af09f7
29861c53
09c31bf3
201c16c3
aabc05dc
2a3c0a57
301c0787
311c1070
ec0c0000
4c8c6b80
00066cac
09c30037
c0bc16c3
09c30a57
24c316c3
0a57f8bc
20261893
183334cd
54cd4006
009017d3
4d6c38c3
ff20323c
716f48c3
61c570cc
62c370cf
763ce04c
72c3f87e
173c206c
12c3fa7e
952b746c
822c333c
fc7e313c
748c42c3
800c233c
fe7e243c
00a7000c
00c70354
323c0494
01938065
049400e7
8035251c
08c30173
608761ec
32c30594
700f6b72
251c0093
500f86dd
323c580c
3203818c
418c223c
ffff001c
ff00011c
68323083
780f3203
323c5c0c
3203818c
418c223c
68323083
7c0f3203
323c440c
3203818c
418c223c
68323083
640f3203
323c500c
3203818c
418c223c
68323083
700f3203
18c309c3
e0bc2ac3
0ab30a40
07875a3c
24c38680
68cc2006
17946007
600768ec
313c1494
404c0030
3f9d243c
180c213c
1070301c
0000311c
6a008c0c
e06c6e80
2187ecef
00b33894
41052025
e4942187
04f382e6
07876a3c
a04c8700
200624c3
35e468cc
68ec1994
87c3e06c
149438e4
0030313c
243c4006
213c3f9d
301c180c
311c1070
8c0c0000
6f006a00
ecefe006
11942187
202500b3
21874105
82c6e294
0133802f
79c360ac
2571775c
0073ec0f
202f2886
e0760296
08040f56
3f36f016
80c3c696
1104301c
0000311c
b05c2c10
605c1b64
a01c1b44
dac30000
106cc01c
0000c11c
0004fe9c
0201065c
065c10c3
303c0209
165c40ac
313c0211
265c81ac
323c0219
6087c1ac
000829dc
0241065c
065c10c3
303c0249
165c40ac
313c0251
465c81ac
243c0259
065cc1ac
10c30261
0269065c
40ac303c
0271165c
81ac313c
0279465c
c1ac343c
219423e4
03e1165c
165c21c3
313c03e9
265c412c
323c03f1
465c81ac
243c03f9
065cc1ac
10c303c1
03c9065c
40ac303c
03d1165c
81ac313c
03d9465c
c1ac343c
413423e4
0281165c
165c21c3
313c0289
265c412c
323c0291
465c81ac
343c0299
39e4c1ac
165c14b4
21c30221
0229165c
412c313c
0231265c
81ac323c
465c06c3
143c0239
d6bcc1ac
03b30a0c
6db739a4
06c11f5c
0285165c
420b333c
4f5c6d77
465c06a1
0d97028d
440b103c
1f5c2d37
165c0681
4d970295
4cf75832
06613f5c
029d365c
0621465c
465c04c3
343c0629
065c402c
303c0631
165c81ac
313c0639
6007c1ac
004492dc
1f3539e4
6cb739a4
06410f5c
0625065c
420b233c
3f5c4c77
365c0621
8c97062d
440b043c
0f5c0c37
065c0601
2c970635
2bf73832
05e12f5c
063d265c
0004299c
0661465c
465c04c3
343c0669
065c402c
303c0671
265c81ac
123c0679
465cc1ac
04c30681
0689465c
402c343c
0691065c
81ac303c
0699265c
c1ac323c
061413e4
16bc06c3
049c0a13
065c0004
20c30201
0209065c
412c303c
0211265c
81ac323c
0219465c
c1ac243c
ffd0323c
6fb46027
0010313c
4f5c6df7
465c06e1
133c0665
2bb7420b
05c12f5c
066d265c
440b433c
0f5c8b77
065c05a1
2dd70675
2b373832
05812f5c
067d265c
0641465c
465c04c3
343c0649
065c402c
303c0651
165c81ac
213c0659
465cc1ac
04c306a1
06a9465c
402c343c
06b1065c
81ac303c
06b9165c
c1ac313c
343c8dd7
123c328d
2af7300d
05612f5c
0625265c
420b413c
0f5c8ab7
065c0541
213c062d
4a77440b
05213f5c
0635365c
98328ad7
0f5c8a37
065c0501
165c063d
21c30221
0229165c
412c313c
0231265c
81ac323c
0239465c
c1ac343c
133c06c3
b0bcfff0
70530a2c
05e1065c
065c40c3
303c05e9
465c422c
343c05f1
065c81ac
303c05f9
6007c1ac
465c1394
04c302e1
02e9465c
402c343c
02f1065c
81ac303c
02f9465c
c1ac343c
d4dc6007
065c002e
20c302e1
02e9065c
412c303c
02f1265c
81ac323c
02f9465c
c1ac343c
0010213c
600740f7
001222dc
00613f5c
0665365c
420b023c
1f5c09f7
165c04e1
323c066d
69b7440b
04c14f5c
0675465c
183200d7
1f5c0977
165c04a1
265c067d
42c30321
0329265c
422c323c
0331465c
81ac343c
0339065c
c1ac303c
088c233c
0161165c
165c41c3
313c0169
465c422c
343c0171
065c81ac
303c0179
433cc1ac
8e77080c
023442e4
1f5c4e77
165c0721
4e5701e5
420b323c
3f5c6937
365c0481
8e5701ed
440b043c
0f5c08f7
065c0461
2e5701f5
28b73832
04412f5c
01fd265c
0161465c
465c04c3
343c0169
065c402c
303c0171
165c81ac
213c0179
4877c1ac
04212f5c
0305265c
433c6857
8837420b
04014f5c
030d465c
103c0857
27f7440b
03e11f5c
0315165c
58324857
3f5c47b7
365c03c1
465c031d
04c30381
0389465c
402c343c
0391065c
81ac303c
0399165c
c1ac313c
2b946027
62126857
6e008857
6c000e57
1f5c6777
165c03a1
333c0305
6737420b
03814f5c
030d465c
103c0757
26f7440b
03611f5c
0315165c
58324757
3f5c46b7
365c0341
8006031d
0385465c
038d465c
0395465c
039d465c
0641065c
065c10c3
303c0649
165c40ac
313c0651
265c81ac
123c0659
465cc1ac
04c306a1
06a9465c
402c343c
06b1065c
81ac303c
06b9465c
c1ac243c
0661065c
065c40c3
303c0669
465c422c
343c0671
065c81ac
303c0679
323cc1ac
413c328d
8677300d
03210f5c
0625065c
420b243c
3f5c4637
365c0301
043c062d
05f7440b
02e11f5c
0635165c
58324657
3f5c45b7
365c02c1
465c063d
04c305e1
05e9465c
402c343c
05f1065c
81ac303c
05f9165c
c1ac713c
680c2cc3
60076c6c
0fb37c94
00613f5c
0665365c
043c80d7
0577420b
02a10f5c
066d065c
213c20d7
4537440b
02812f5c
0675265c
783260d7
4f5c64f7
465c0261
065c067d
10c30641
0649065c
40ac303c
0651165c
81ac313c
0659465c
c1ac243c
06a1065c
065c10c3
303c06a9
165c40ac
313c06b1
465c81ac
343c06b9
00d7c1ac
328d303c
300d423c
0f5c84b7
065c0241
243c0625
4477420b
02213f5c
062d365c
440b043c
1f5c0437
165c0201
44970635
43f75832
01e13f5c
063d365c
0221465c
465c04c3
343c0229
065c402c
303c0231
06c381ac
0239265c
c1ac123c
0a0cd6bc
0861465c
465c04c3
343c0869
065c402c
303c0871
165c81ac
613c0879
37f3c1ac
366407c3
201c7c2c
211cdddd
42c3dddd
64dc34e4
065c001a
10c30481
0489065c
40ac303c
0491165c
81ac313c
0499265c
c1ac323c
0010033c
1f5c03b7
165c01c1
303c0485
6377420b
01a14f5c
048d465c
440b103c
2f5c2337
265c0181
63970495
62f77832
01614f5c
049d465c
1c2f0006
21c33a89
313c3aa9
5ac9412c
81ac323c
343c9ae9
6087c1ac
7def5194
640c1cc3
64d26ccc
366407c3
2ac3a0c3
02dc4007
9b090016
9b2904c3
402c343c
303c1b49
3b6981ac
c1ac213c
04e1465c
465c04c3
343c04e9
065c402c
303c04f1
165c81ac
413c04f9
065cc1ac
10c30501
0509065c
40ac303c
0511165c
81ac313c
0519065c
c1ac303c
20066037
0006111c
065c2077
10c30521
0529065c
40ac303c
0531165c
81ac313c
0539065c
c1ac303c
08c360b7
34c317c3
0a22a0bc
20c62373
5b093def
5b2942c3
422c323c
343c9b49
1b6981ac
c1ac303c
3b897e0f
3ba921c3
412c313c
323c5bc9
9be981ac
c1ac343c
065c7e2f
10c30101
0109065c
40ac303c
0111165c
81ac313c
0119265c
c1ac323c
465c7e4f
04c30121
0129465c
402c343c
0131065c
81ac303c
0139165c
c1ac313c
265c7e6f
42c30a21
0a29265c
422c323c
0a31465c
81ac343c
0a39065c
c1ac303c
3e8f2c4c
0a21265c
265c42c3
323c0a29
465c422c
343c0a31
065c81ac
303c0a39
2c6cc1ac
265c3eaf
42c30a21
0a29265c
422c323c
0a31465c
81ac343c
0a39065c
c1ac303c
3ecf2c8c
0a21265c
265c42c3
323c0a29
465c422c
343c0a31
065c81ac
303c0a39
2cacc1ac
265c3eef
42c30a21
0a29265c
422c323c
0a31465c
81ac343c
0a39065c
c1ac303c
1cc37f0f
6ccc640c
07c364d2
d0c33664
40072dc3
000832dc
700c4cc3
08c3bccc
31a4005c
8e4c0037
17c308c3
35c340c6
0e934664
055440e7
03544127
6e944167
0010313c
4f5c6e37
465c0701
133c0665
22b7420b
01412f5c
066d265c
440b433c
0f5c8277
065c0121
2e170675
22373832
01012f5c
067d265c
0641465c
465c04c3
343c0649
065c402c
303c0651
165c81ac
213c0659
465cc1ac
04c306a1
06a9465c
402c343c
06b1065c
81ac303c
06b9165c
c1ac313c
343c8e17
123c328d
21f7300d
00e12f5c
0625265c
420b413c
0f5c81b7
065c00c1
213c062d
4177440b
00a13f5c
0635365c
983281d7
0f5c8137
065c0081
165c063d
21c30221
0229165c
412c313c
0231265c
81ac323c
0239465c
c1ac343c
133c06c3
12bcfff0
065c0a58
10c30861
0869065c
40ac303c
0871165c
81ac313c
0879265c
c1ac623c
ffffb21c
60073bc3
ffb024dc
fc763a96
08040f56
3f36f016
40c3c596
301c81c3
311c1110
6c0c0000
eebc2c10
50c309f8
08c35264
2006606c
0002111c
60073183
245c1354
02c30221
0229245c
402c323c
0231045c
81ac303c
245c04c3
123c0239
d6bcc1ac
08c30a0c
2006606c
0010111c
60073183
005fd2dc
0201245c
245c02c3
323c0209
045c402c
303c0211
145c81ac
313c0219
60a7c1ac
000804dc
0a01045c
045c10c3
303c0a09
145c40ac
313c0a11
245c81ac
323c0a19
6007c1ac
a0076e54
09c31f54
05d9305c
1a1435e4
03c7353c
6d00402c
6e376d8b
12546007
07013f5c
06c5345c
08320e17
1f5c0df7
145c06e1
400606cd
06d5245c
06dd245c
301c03d3
311c106c
6c0c0000
0ca96c0c
0cc910c3
40ac103c
2db701c3
06c11f5c
06c5145c
483220c3
3f5c4d77
345c06a1
000606cd
06d5045c
06dd045c
145c2006
145c06e5
145c06ed
145c06f5
245c06fd
02c30241
0249245c
402c323c
0251045c
81ac303c
0259145c
c1ac313c
fff0233c
602c08c3
139432e4
0221245c
245c02c3
323c0229
045c402c
303c0231
04c381ac
0239245c
c1ac123c
0a0cd6bc
ec4c38c3
0221045c
045c10c3
303c0229
145c40ac
313c0231
245c81ac
323c0239
73e4c1ac
145c3594
21c305c1
05c9145c
412c313c
05d1245c
81ac323c
05d9045c
c1aca03c
0601145c
145c21c3
313c0609
245c412c
323c0611
045c81ac
903c0619
18c3c1ac
2d37246c
06812f5c
02e5245c
ffff141c
28322d37
0f5c2cf7
045c0661
200602ed
02f5145c
02fd145c
245c4093
02c305e1
05e9245c
402c323c
05f1045c
81ac303c
05f9145c
c1ac613c
106c301c
0000311c
6c6c6c0c
06c363d2
c0073664
001382dc
201c782c
211cdddd
02c3dddd
14dc30e4
796c0014
323c4c2c
3203818c
418c223c
ffff101c
ff00111c
533c3183
5203408c
684c28c3
04dc35e4
145c000f
21c30361
0369145c
412c313c
0371245c
81ac323c
0379045c
c1ac103c
2ef22cb7
145c2026
2f5c0365
245c0641
32c3036d
0375345c
045c02c3
145c037d
21c30361
0369145c
412c313c
0371245c
81ac323c
0379045c
c1ac303c
0010233c
3f5c4e77
345c0721
123c0365
2c77420b
06212f5c
036d245c
033c6e57
0c37440b
06010f5c
0375045c
38322e57
2f5c2bf7
245c05e1
6e57037d
008703c3
145c3c35
21c30161
0169145c
412c313c
0171245c
81ac323c
0179045c
c1ac203c
0301145c
145c01c3
313c0309
045c402c
303c0311
145c81ac
313c0319
6980c1ac
2f5c6bb7
245c05c1
033c0305
0b77420b
05a11f5c
030d145c
323c4b97
6b37440b
05813f5c
0315345c
18320b97
1f5c0af7
145c0561
02f3031d
32c34e57
13946087
045c0026
20060625
062d145c
0635145c
063d145c
0385045c
038d145c
0395145c
039d145c
0621245c
245c02c3
323c0629
045c402c
303c0631
145c81ac
213c0639
4007c1ac
045c3f54
10c30661
0669045c
40ac303c
0671145c
81ac313c
0679045c
c1ac303c
2e946007
0010323c
088c233c
0f5c4eb7
045c0741
233c0625
4ab7424b
05410f5c
062d045c
444b233c
0f5c4a77
045c0521
233c0635
4a37c88c
05013f5c
063d345c
0ef20e97
145c2026
2f5c0625
245c0741
32c3062d
0635345c
045c02c3
145c063d
21c30361
0369145c
412c313c
0371245c
81ac323c
0379045c
c1ac303c
05946087
084c29c3
0a64e6bc
0221045c
045c10c3
303c0229
145c40ac
313c0231
245c81ac
723c0239
b01cc1ac
75e40000
b01c1bb4
03130001
0221045c
045c10c3
303c0229
145c40ac
313c0231
245c81ac
523c0239
75c3c1ac
00d3b6c3
ac2c38c3
b01c75c3
045c0000
10c30241
0249045c
40ac303c
0251145c
81ac313c
0259045c
c1ac203c
642c18c3
159432e4
29f7246c
04e12f5c
02e5245c
ffff141c
283229f7
0f5c29b7
045c04c1
200602ed
02f5145c
02fd145c
0000901c
c01ca9c3
c11c106c
0d730000
680c2cc3
63d26c6c
366406c3
001c782c
011cdddd
10c3dddd
5f9431e4
686c596c
818c133c
033c1303
482c418c
818c323c
d23c3203
201c418c
211cffff
3283ff00
3d036832
58ccd3c3
301cd284
311cffff
1383ff00
408c313c
7c323003
0dc36212
1bc341a0
08c328f2
32e4604c
37e43614
06730d35
604c08c3
043425e4
041435e4
35e40593
32e40314
28c32814
4977486c
04a13f5c
02e5345c
ffff241c
48324977
1f5c4937
145c0481
400602ed
02f5245c
02fd245c
32c3584c
eeee001c
eeee011c
333c3003
33c40b0d
a21c7f52
96c30001
638362c3
9594c007
20071ac3
28c33194
045c284c
20c30221
0229045c
412c303c
0231245c
81ac323c
0239045c
c1ac203c
0b5412e4
600767a0
003097dc
12c304c3
0a0cd6bc
60730ac3
03c1245c
245c02c3
323c03c9
045c402c
303c03d1
245c81ac
323c03d9
64f2c1ac
d6bc04c3
045c0a0c
10c30361
0369045c
40ac303c
0371145c
81ac313c
0379245c
c1ac323c
53546007
1e353ae4
68f73aa4
04612f5c
0365245c
420b033c
1f5c08b7
145c0441
48d7036d
440b323c
3f5c6877
345c0421
08d70375
08371832
04011f5c
037d145c
40060693
0365245c
036d245c
0375245c
037d245c
01e1045c
045c10c3
303c01e9
145c40ac
313c01f1
245c81ac
023c01f9
07f7c1ac
03e13f5c
0305345c
420b103c
2f5c27b7
245c03c1
67d7030d
440b033c
0f5c0777
045c03a1
27d70315
27373832
03812f5c
031d245c
0301045c
045c10c3
303c0309
145c40ac
313c0311
045c81ac
203c0319
145cc1ac
01c301e1
01e9145c
402c313c
01f1045c
81ac303c
01f9145c
c1ac313c
313523e4
01c1145c
145c01c3
313c01c9
045c402c
303c01d1
145c81ac
313c01d9
141dc1ac
62f23320
6d006026
2f5c66f7
245c0361
033c0305
06b7420b
03411f5c
030d145c
323c46d7
6677440b
03213f5c
0315345c
183206d7
1f5c0637
145c0301
0593031d
0161045c
045c10c3
303c0169
145c40ac
313c0171
045c81ac
303c0179
6d00c1ac
1f5c65f7
145c02e1
333c0305
65b7420b
02c10f5c
030d045c
213c25d7
4577440b
02a12f5c
0315245c
783265d7
0f5c6537
045c0281
145c031d
21c302e1
02e9145c
412c313c
02f1245c
81ac323c
02f9045c
c1ac103c
145c24f7
21c30301
0309145c
412c313c
0311245c
81ac323c
0319045c
c1ac303c
21c324d7
1b3532e4
02613f5c
0305345c
420b113c
1f5c24b7
145c0241
44d7030d
440b323c
3f5c6477
345c0221
04d70315
04371832
02011f5c
031d145c
40072ac3
001d12dc
09a1045c
045c10c3
303c09a9
145c40ac
313c09b1
245c81ac
523c09b9
a007c1ac
045c2754
10c305c1
05c9045c
40ac303c
05d1145c
81ac313c
05d9245c
c1ac123c
05a1045c
045c20c3
303c05a9
245c412c
323c05b1
045c81ac
203c05b9
12e4c1ac
0ac30714
32e46420
04c30334
245c5664
02c305e1
05e9245c
402c323c
05f1045c
81ac303c
05f9145c
c1ac613c
0601245c
245c02c3
323c0609
045c402c
303c0611
145c81ac
313c0619
93e4c1ac
39c37054
345c6d09
09c305e5
045c0129
19c305ed
145c2549
29c305f5
245c4969
045c05fd
10c305c1
05c9045c
40ac303c
05d1145c
81ac313c
05d9245c
c1ac323c
63f73aa4
01e11f5c
05c5145c
420b333c
0f5c63b7
045c01c1
23d705cd
440b213c
2f5c4377
245c01a1
63d705d5
63377832
01810f5c
05dd045c
0641145c
145c21c3
313c0649
245c412c
323c0651
045c81ac
103c0659
01c3c1ac
1f5c22f7
145c0161
303c0625
62b7420b
01413f5c
062d345c
440b103c
1f5c2277
145c0121
42d70635
42375832
01013f5c
063d345c
045c0006
045c0665
045c066d
045c0675
0ff3067d
145c2006
145c05e5
145c05ed
145c05f5
145c05fd
145c0605
145c060d
145c0615
145c061d
145c05c5
145c05cd
145c05d5
245c05dd
02c30201
0209245c
402c323c
0211045c
81ac303c
0219145c
c1ac313c
055460e7
03546127
35946167
0641245c
245c02c3
323c0649
045c402c
303c0651
145c81ac
213c0659
12c3c1ac
2f5c41f7
245c00e1
013c0625
01b7420b
00c10f5c
062d045c
440b213c
2f5c4177
245c00a1
61d70635
61377832
00810f5c
063d045c
145c2006
145c0665
145c066d
145c0675
03b3067d
02e1245c
245c02c3
323c02e9
045c402c
303c02f1
145c81ac
313c02f9
6dd2c1ac
245c4006
245c0625
245c062d
245c0635
0073063d
00b367c3
106c801c
0000811c
301cf84c
311caaaa
784faaaa
fbc4265c
600c08c3
2f696c0c
09692cd2
341c30c3
6cf20004
dddd101c
dddd111c
00d3382f
dddd201c
dddd211c
782c582f
dddd001c
dddd011c
31e410c3
796c5d94
323c4c6c
3203818c
418c223c
ffff001c
ff00011c
68323083
7c323203
100c533c
0321145c
145c21c3
313c0329
245c412c
323c0331
045c81ac
103c0339
58ccc1ac
13e46aa0
65201f35
60f76e80
00611f5c
0325145c
420b333c
0f5c60b7
045c0041
20d7032d
440b213c
2f5c4077
245c0021
60d70335
60377832
00010f5c
033d045c
20060153
0325145c
032d145c
0335145c
033d145c
680c28c3
4bd24d2c
0a41045c
341c30c3
65d20001
04c378cc
26642ea0
66bc06c3
a21c0a40
1ac3ffff
54dc2007
0026fff7
fc763b96
08040f56
fc967016
105c40c3
21c305e1
05e9105c
412c313c
05f1205c
81ac323c
05f9105c
c1ac013c
245c4006
245c05e5
245c05ed
245c05f5
245c05fd
245c0605
245c060d
245c0615
6e24061d
4004633c
f5240733
301ca04c
311caaaa
604faaaa
f324c2d2
0a4066bc
05c1145c
145c21c3
313c05c9
245c412c
323c05d1
145c81ac
313c05d9
133cc1ac
20f7fff0
00612f5c
05c5245c
420b113c
2f5c20b7
245c0041
60d705cd
440b133c
1f5c2077
145c0021
40d705d5
40375832
00013f5c
05dd345c
145c05c3
21c305c1
05c9145c
412c313c
05d1245c
81ac323c
05d9145c
c1ac313c
b8946007
0e560496
00000804
0136f016
61c350c3
83c372c3
106c301c
0000311c
6d4c6c0c
12c367d2
366426c3
600730c3
40066b54
2e24580f
744cf524
21546007
744f7fe5
4c6c74ec
400654ef
4c2f4c6f
4ccf4c8f
4b804d2c
4d8f4d6f
4cef4006
201c4d0f
211caaaa
4c4faaaa
235c4006
408601c5
40064def
780f4f0f
081302c3
6025748c
0026748f
600738c3
74ac3954
74af6c00
11b4301c
0000311c
201c8c0c
211cb638
534f0014
d3efb36f
756cf3cf
738f6bd2
4fac756c
756c53af
8f8f6fac
8faf756c
956f0093
93af938f
6025758c
6186758f
4026718f
201c51cf
211c1250
680c0000
680f6025
313c1271
62d24004
04c3f324
09f1a4bc
0424045c
313c00b3
62d24004
8076f324
08040f56
0136f016
60c3ff96
72c341c3
9abc83c3
5f3c0bae
053c0040
06c3fe7e
2fc314c3
0bae9ebc
1d740007
0100463c
9abc04c3
00370bae
17c304c3
9ebc2fc3
00070bae
463c1074
04c30200
0bae9abc
04c30037
2fc318c3
0bae9ebc
000630c3
021530e4
01961fe6
0f568076
00000804
ff967016
41c360c3
0bae9abc
100f0037
1110301c
0000311c
335c6c0c
36640784
1fe650c3
3354a007
15c306c3
9ebc2fc3
00070bae
05c32074
d4a8101c
0014111c
eabc4017
802608cb
17540007
101c05c3
111cd4c0
40170014
08cbeabc
0dd28046
101c05c3
111cd4dc
40170014
08cbeabc
03d28086
00ff401c
1110301c
0000311c
335c6c0c
05c307c4
04c33664
0e560196
00000804
60c3f016
73c352c3
24c38157
0bae92bc
13740007
0100063c
24c315c3
0bae92bc
0b740007
0200063c
24c317c3
0bae92bc
000630c3
021530e4
0f561fe6
00000804
0336f016
80c3fd96
00c02f3c
023c0006
901cfe7e
911c10f8
09c30000
6d4c600c
12c301c3
00773664
1110401c
0000411c
335c700c
00970784
50c33664
335c700c
00970784
60c33664
335c700c
00970784
70c33664
3b54a007
3954c007
37540007
15c308c3
37c326c3
0a4edabc
2f740007
209705c3
0a7352bc
209706c3
0a7352bc
209707c3
0a7352bc
600c09c3
2f5c8e6c
02c30021
26c315c3
466437c3
209705c3
0a7352bc
209706c3
0a7352bc
209707c3
0a7352bc
60376097
15c308c3
37c326c3
0a4f5abc
800630c3
021534e4
aad29fe6
1110301c
0000311c
335c6c0c
05c307c4
cad23664
1110301c
0000311c
335c6c0c
06c307c4
ead23664
1110301c
0000311c
335c6c0c
07c307c4
04c33664
c0760396
08040f56
3f36f016
b0c3fa96
1f3cd1c3
00060180
fe7e013c
10f8c01c
0000c11c
600c0cc3
02c36d4c
01373664
1110401c
0000411c
335c700c
01570784
50c33664
335c700c
01570784
60c33664
335c700c
01570784
70c33664
335c700c
01570784
80c33664
335c700c
01570784
90c33664
335c700c
01570784
a0c33664
4d54a007
4b54c007
4954e007
400728c3
39c34654
43546007
41540007
15c30bc3
37c326c3
0a4edabc
600730c3
05c33874
52bc2157
06c30a73
52bc2157
07c30a73
52bc2157
2cc30a73
0006680c
00050f5c
00278f5c
00479f5c
0067af5c
2f5c8e4c
02c30081
26c315c3
466437c3
215708c3
0a7352bc
215709c3
0a7352bc
21570ac3
0a7352bc
60376157
18c30dc3
3ac329c3
0a4f5abc
800630c3
021534e4
aad29fe6
1110301c
0000311c
335c6c0c
05c307c4
cad23664
1110301c
0000311c
335c6c0c
06c307c4
ead23664
1110301c
0000311c
335c6c0c
07c307c4
28c33664
301c4ad2
311c1110
6c0c0000
07c4335c
366408c3
6ad239c3
1110301c
0000311c
335c6c0c
09c307c4
0ac33664
301c09d2
311c1110
6c0c0000
07c4335c
04c33664
fc760696
08040f56
3f36f016
0337f196
42b722f7
03c01f3c
213c4006
201cfe7e
211c10f8
480c0000
03c3494c
03772664
1110401c
0000411c
335c700c
03970784
50c33664
335c700c
03970784
60c33664
335c700c
03970784
70c33664
335c700c
03970784
80c33664
335c700c
03970784
90c33664
335c700c
03970784
a0c33664
335c700c
03970784
b0c33664
335c700c
03970784
c0c33664
335c700c
03970784
d0c33664
7654a007
7454c007
7254e007
600738c3
29c36f54
6c544007
60073ac3
2bc36954
66544007
60073cc3
00076354
03176154
26c315c3
dabc37c3
00070a4e
02d75974
29c318c3
dabc3ac3
00070a4e
05c35174
52bc2397
06c30a73
52bc2397
07c30a73
52bc2397
08c30a73
52bc2397
09c30a73
52bc2397
0ac30a73
52bc2397
301c0a73
311c10f8
6c0c0000
8f5ce037
9f5c0027
af5c0047
40060067
00852f5c
00a52f5c
00c52f5c
00e7bf5c
0107cf5c
0127df5c
3f5c8e2c
03c301a1
25c312c3
466436c3
23970bc3
0a7352bc
23970cc3
0a7352bc
23970dc3
0a7352bc
40374397
1bc30297
3dc32cc3
0a4f5abc
04e48006
9fe60215
301caad2
311c1110
6c0c0000
07c4335c
366405c3
301ccad2
311c1110
6c0c0000
07c4335c
366406c3
301cead2
311c1110
6c0c0000
07c4335c
366407c3
6ad238c3
1110301c
0000311c
335c6c0c
08c307c4
29c33664
301c4ad2
311c1110
6c0c0000
07c4335c
366409c3
6ad23ac3
1110301c
0000311c
335c6c0c
0ac307c4
2bc33664
301c4ad2
311c1110
6c0c0000
07c4335c
36640bc3
6ad23cc3
1110301c
0000311c
335c6c0c
0cc307c4
2dc33664
301c4ad2
311c1110
6c0c0000
07c4335c
36640dc3
0f9604c3
0f56fc76
00000804
3f36f016
d0c3f396
427722b7
03406f3c
263c4006
201cfe7e
211c10f8
480c0000
03c3494c
266416c3
401c02f7
411c1110
700c0000
0784335c
36640317
700c70c3
0784335c
36640317
700c80c3
0784335c
36640317
700c50c3
0784335c
36640317
700c90c3
0784335c
36640317
700ca0c3
0784335c
36640317
700cb0c3
0784335c
36640317
e007c0c3
38c37654
73546007
7154a007
400729c3
3ac36e54
6b546007
40072bc3
00076854
02976654
28c317c3
dabc35c3
00070a4e
0dc35e74
0bae9abc
0dc30337
26c319c3
0bae9ebc
53740007
231709c3
0a7352bc
231707c3
0a7352bc
231708c3
0a7352bc
101c05c3
111cd4fc
43170014
08cbeabc
05c305d2
52bc2317
301c0a73
311c10f8
6c0c0000
8f5ce037
a0b70027
2f5c4006
2f5c0065
2f5c0301
40060085
00a52f5c
00c7af5c
00e7bf5c
0107cf5c
3f5c8e0c
03c30161
39c312c3
0ac34664
52bc2317
0bc30a73
52bc2317
46170a73
0cc345f2
52bc2317
63170a73
02576037
2bc31ac3
5abc3cc3
80060a4f
021504e4
ead29fe6
1110301c
0000311c
335c6c0c
07c307c4
38c33664
301c6ad2
311c1110
6c0c0000
07c4335c
366408c3
301caad2
311c1110
6c0c0000
07c4335c
366405c3
4ad229c3
1110301c
0000311c
335c6c0c
09c307c4
3ac33664
301c6ad2
311c1110
6c0c0000
07c4335c
36640ac3
4ad22bc3
1110301c
0000311c
335c6c0c
0bc307c4
3cc33664
301c6ad2
311c1110
6c0c0000
07c4335c
36640cc3
0d9604c3
0f56fc76
00000804
0bfb0cbc
00000804
0bfafcbc
00000804
0bfb26bc
00000804
1f36f016
b1c350c3
c2c3b264
400cc264
1110301c
0000311c
640c2c0c
04c38c6c
385420e4
36544047
f680853c
07a4315c
366414cc
901c60c3
911c0ef0
a01c0000
a11c0bb4
753c0000
0007f6c0
49c31194
1ac3700c
17c3040c
301c3664
311c0b84
6c0c0000
2227001c
00263664
301c07d3
311c1118
6c0c0000
08c38d4c
2bc316c3
4664758b
680c29c3
100c4ac3
366417c3
d56c0053
1118301c
0000311c
440c2c0c
03c73c3c
6c00082c
0c6c856c
54cc16c3
356c4664
62e421c3
301c0a54
311c1110
6c0c0000
07c4335c
01b306c3
66bc05c3
30c30a40
301c6ad2
311c0b84
6c0c0000
2225001c
00063664
0f56f876
00000804
3f36f016
a1c3fb96
0264d3c3
c264c2c3
41374006
301c40f7
311c1110
6c0c0000
303c2c10
83c303c7
302c49c3
18c38184
e007e46c
000c52dc
1e79375c
09dc6127
203c000c
303cfff0
7fe500b6
b33c32a3
3bc3f88c
644c67f2
18546007
80078c89
301c1594
311c1118
4c0c0000
1388301c
0000311c
a112ac0b
01003f3c
898c6037
1f3c07c3
25c300c0
18c302b3
62c34749
0001641c
1118501c
0000511c
00c01f3c
01000f3c
740cc9d2
51cb48c3
8d8c0037
600607c3
740c0113
8d8c0037
201c07c3
36c305b4
60c34664
00d6001c
febd631c
001c7854
631c00d5
7354feab
7074c007
88f24bc3
644c18c3
2c546007
40074c89
301c2994
311c1388
6c0b0000
63e46112
19c31bd4
1ac3046c
3dc34006
0a4e5abc
12940007
680c2ac3
846c19c3
03c30037
26c320d7
6ebc34c3
00070a0a
2ac33f54
66bc080c
301c0a40
311c1118
6c0c0000
66c60593
c31c60b7
03540004
20b72946
0bb4301c
0000311c
6c2c6c0c
6c2b6c0c
1118501c
0000511c
08b46027
6dac740c
366407c3
00d5001c
740c0493
80378006
00411f5c
00251f5c
00068dcc
20c316c3
466460d7
740c06f2
07c36dac
02133664
0580303c
680f2ac3
301cc38f
311c1118
6c0c0000
07c36dac
00063664
00260053
fc760596
08040f56
fb967016
61c330c3
326452c3
301c6137
311c1118
6c0c0000
301c8c2c
311c1179
2f5c0000
4c0d0081
68d2700c
2abc04c3
04c309df
9cbc2586
301c08cb
311c1118
6c0c0000
201c6d2c
403700c8
40264077
458640b7
04c340f7
d51c101c
0014111c
611723c3
09dea8bc
05c3c5d2
0ba2d8bc
05c30093
0ba1a6bc
002710c3
05c30b54
0b9ffabc
ffe0303c
31e42026
101c0335
01c300d2
0e560596
00000804
f6963016
046c40c3
400630c3
0010211c
60073283
000b62dc
0221545c
545c25c3
353c0229
245c412c
323c0231
545c81ac
253c0239
644cc1ac
34dc32e4
4006000a
0001211c
02770283
1a940007
345c6106
5f5c0205
545c0121
15c3020d
0215145c
245c25c3
35c3021d
0625345c
062d545c
145c15c3
25c30635
063d245c
b1091c73
b12915c3
40ac353c
313c3149
516981ac
c1ac523c
aad2a237
345c6026
a0060205
020d545c
0215545c
20460193
0205145c
01012f5c
020d245c
345c32c3
52c30215
021d545c
145c2006
145c0625
145c062d
145c0635
245c063d
52c30241
0249245c
42ac323c
0251545c
81ac353c
0259145c
c1ac313c
0010533c
1f5ca1f7
145c00e1
353c0245
61b7420b
00c15f5c
024d545c
213c21d7
4177440b
00a12f5c
0255245c
783261d7
5f5c6137
545c0081
145c025d
21c30221
0229145c
412c313c
0231245c
81ac323c
545c04c3
153c0239
d6bcc1ac
145c0a0c
21c30801
0809145c
412c313c
0811245c
81ac323c
0819545c
c1ac353c
68546007
1000043c
38bc2006
0c530a57
200630c3
0001111c
60073183
41265b54
0205245c
345c6006
345c020d
345c0215
545c021d
15c30241
0249545c
40ac353c
0251145c
81ac313c
0259245c
c1ac323c
0010133c
2f5c20f7
245c0061
513c0245
a0b7420b
00411f5c
024d145c
323c40d7
6077440b
00213f5c
0255345c
b832a0d7
1f5ca037
145c0001
245c025d
52c30221
0229245c
42ac323c
0231545c
81ac353c
245c04c3
123c0239
d6bcc1ac
545c0a0c
15c30941
0949545c
40ac353c
0951145c
81ac313c
0959245c
c1ac323c
04c363d2
545c3664
15c30201
0209545c
40ac353c
0211145c
81ac313c
0219245c
c1ac323c
60277fe5
145c24b4
21c30921
0929145c
412c313c
0931245c
81ac323c
0939545c
c1ac353c
11946007
0901145c
145c21c3
313c0909
245c412c
323c0911
545c81ac
353c0919
63d2c1ac
366404c3
0c560a96
00000804
fb961016
646c40c3
111c2006
31830001
82dc6007
4109000b
412912c3
40ac323c
313c2149
416981ac
c1ac123c
2cd22137
305c6026
20060205
020d105c
0215105c
021d105c
404601d3
0205205c
00813f5c
020d305c
105c13c3
23c30215
021d205c
345c6006
345c0625
345c062d
345c0635
145c063d
21c30241
0249145c
412c313c
0251245c
81ac323c
0259145c
c1ac313c
0010133c
2f5c20f7
245c0061
113c0245
20b7420b
00412f5c
024d245c
133c60d7
2077440b
00211f5c
0255145c
583240d7
3f5c4037
345c0001
145c025d
21c30221
0229145c
412c313c
0231245c
81ac323c
245c04c3
123c0239
d6bcc1ac
145c0a0c
21c30801
0809145c
412c313c
0811245c
81ac323c
0819145c
c1ac313c
043c66d2
20061000
0a5738bc
0941245c
245c12c3
323c0949
145c40ac
313c0951
245c81ac
323c0959
63d2c1ac
366404c3
0921145c
145c21c3
313c0929
245c412c
323c0931
145c81ac
313c0939
6007c1ac
245c1194
12c30901
0909245c
40ac323c
0911145c
81ac313c
0919245c
c1ac323c
04c363d2
05963664
08040856
0f36f016
41c350c3
002672c3
e000011c
41e410c3
655c2054
301c13e4
311c106c
6c0c0000
b35c6c0c
40060079
a23c0213
363c100c
34e42a1d
955c0994
09c31404
60811ac3
78e483c3
40250654
f0142be4
00530006
f0760026
08040f56
f5244e24
2464305c
323c69f2
62d24004
01c3f324
0a4066bc
305c03d3
241c2484
6cd20400
24a4305c
60062c2f
105c642f
400724a7
f3241054
105c01d3
105c2487
642f24a7
f32442d2
01fc021c
40062406
09e0bebc
00000804
20c33016
2e2441c3
000cf524
1f540007
03e4638c
60060494
00f3680f
438c680f
abafa3ac
4f8f63ac
634f6006
1250201c
0000211c
6025680c
313c680f
62d24004
405cf324
02bc0427
00b309f1
4004313c
f32462d2
08040c56
50c33016
1074401c
0000411c
3fe604c3
09e2f6bc
752f6006
76bc04c3
0c5609e4
00000804
63c3f016
f524ae24
11b4301c
0000311c
600c8c0c
738f6bd2
efac600c
600cf3af
8f8f6fac
8faf600c
800f0093
93af938f
536f334f
718f6186
f1cfe026
1250201c
0000211c
6f80680c
6157680f
353c726f
62d24004
06c3f324
09e476bc
a4bc04c3
0f5609f1
00000804
50c3f016
72c361c3
0e00403c
3fe604c3
09e2f6bc
0447363c
735c7580
04c32667
09e476bc
0f560006
00000804
0336f016
40c3f896
82c371c3
a3d793c3
0e00603c
3fe606c3
09e2f6bc
1494a027
00478f5c
00679f5c
628681b7
273c6037
323c0447
71804a80
710061f7
2744335c
36640fc3
a3d20053
68f26057
0447373c
835c7180
935c25a7
06c325c7
09e476bc
a0270006
00570294
c0760896
08040f56
ff967016
61c350c3
403c4037
04c30e00
f6bc3fe6
363c09e2
75800447
00012f5c
256d235c
76bc04c3
000609e4
0e560196
00000804
0136f016
50c3f496
005c71c3
10c304c1
04c9055c
40ac303c
04d1155c
81ac313c
04d9255c
c1ac823c
64c39689
343c96a9
d6c9432c
81ac363c
403c16e9
18c3c1ac
06e4015c
02c01f3c
0b948087
60064706
0a4e5abc
54dc0007
62d70024
11f38def
60064706
0a4e5abc
b4dc0007
62d70023
8def80c6
655c42d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8a8f8c4c
655c42d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8aaf8c6c
655c42d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8acf8c8c
655c42d7
06c30a21
0a29655c
402c363c
0a31055c
81ac303c
0a39155c
c1ac313c
8aef8cac
d70942d7
d72906c3
402c363c
303c1749
376981ac
c1ac313c
42d76a0f
64c39789
343c97a9
d7c9432c
81ac363c
303c17e9
6a2fc1ac
155c42d7
41c30101
0109155c
422c313c
0111455c
81ac343c
0119655c
c1ac363c
42d76a4f
0121055c
055c10c3
303c0129
155c40ac
313c0131
455c81ac
343c0139
6a6fc1ac
655c42d7
06c30181
0189655c
402c363c
0191055c
81ac303c
0199155c
c1ac313c
42d768ef
01a1455c
455c64c3
343c01a9
655c432c
363c01b1
055c81ac
303c01b9
690fc1ac
696c42d7
698f6285
228662d7
62d72ccf
7589cd6c
75a943c3
422c233c
0141455c
455c04c3
343c0149
055c402c
303c0151
155c81ac
313c0159
323cc1ac
780f81ac
255cf82f
42c30241
0249255c
422c323c
0251455c
81ac343c
0259055c
c1ac303c
155c784f
21c303c1
03c9155c
412c313c
03d1255c
81ac323c
03d9455c
c1ac343c
011c0006
30a35011
2006786f
255c388f
42c30241
0249255c
422c323c
0251455c
81ac343c
0259055c
c1ac103c
1f5c22b7
155c0141
42970265
420b323c
3f5c6277
355c0121
8297026d
440b043c
0f5c0237
055c0101
22970275
21f73832
00e12f5c
027d255c
03c1455c
455c04c3
343c03c9
055c402c
303c03d1
155c81ac
213c03d9
41b7c1ac
00c12f5c
03e5255c
433c6197
8177420b
00a14f5c
03ed455c
103c0197
2137440b
00811f5c
03f5155c
58324197
3f5c40f7
355c0061
580c03fd
818c323c
223c3203
401c418c
411cffff
3483ff00
32036832
582c780f
818c323c
223c3203
3483418c
32036832
584c782f
818c323c
223c3203
3483418c
32036832
586c784f
818c323c
223c3203
3483418c
32036832
588c786f
818c323c
223c3203
3483418c
32036832
3689788f
36a921c3
412c313c
323c56c9
96e981ac
c1ac343c
13946087
0181155c
155c21c3
313c0189
255c412c
323c0191
455c81ac
343c0199
733cc1ac
02530140
0a21055c
055c10c3
303c0a29
155c40ac
313c0a31
255c81ac
323c0a39
733cc1ac
42d70080
353c88cc
60370180
20c602c3
37c324c3
0a3f38bc
233c30e3
323c800c
3203818c
418c223c
ffff401c
ff00411c
68323483
788f3203
06c3d689
363cd6a9
16c9402c
81ac303c
313c36e9
22d7c1ac
44946087
64c39709
343c9729
d749432c
81ac363c
203c1769
455cc1ac
64c304e1
04e9455c
432c343c
04f1655c
81ac363c
04f9055c
c1ac403c
0501655c
655c06c3
363c0509
055c402c
303c0511
655c81ac
363c0519
6037c1ac
011c0006
00770006
0521655c
655c06c3
363c0529
055c402c
303c0531
655c81ac
363c0539
60b7c1ac
34c308c3
0a22a0bc
055c0453
20c30a21
0a29055c
412c303c
0a31255c
81ac323c
0a39455c
c1ac343c
42d7670f
106c301c
0000311c
a8cc6c0c
665c68c3
c03731a4
08c38e4c
40c612c3
466435c3
80760c96
08040f56
00000804
f8963016
8e24236c
634cf524
62dc6007
20070008
000832dc
52c34409
323c4429
a44942ac
81ac353c
323c4469
501cc1ac
511c5020
25c35544
709432e4
634f6006
a1f7a38c
0a9405e4
02c5315c
02cd315c
02d5315c
02dd315c
5f5c0433
515c00e1
41d702c5
420b323c
3f5c61b7
315c00c1
a1d702cd
440b253c
2f5c4177
215c00a1
61d702d5
61377832
00815f5c
02dd515c
63ac438c
63ac6baf
515c4f8f
25c302e1
02e9515c
412c353c
02f1215c
81ac323c
02f9515c
c1ac353c
fff0533c
2f5ca0f7
215c0061
553c02e5
a0b7420b
00412f5c
02ed215c
533c60d7
a077440b
00215f5c
02f5515c
583240d7
3f5c4037
315c0001
618c02fd
12946187
205c4026
201c0427
211c1250
680c0000
680f6025
4004343c
f32462d2
09f102bc
343c00b3
62d24004
0896f324
08040c56
236c3016
f5248e24
6007634c
20073354
640c3154
434b201c
5041211c
35e452c3
40062994
438c434f
049402e4
a56fa006
656c0153
029430e4
438c456f
6baf63ac
4f8f63ac
7fe5658c
618c658f
12946187
205c4026
201c0427
211c1250
680c0000
680f6025
4004343c
f32462d2
09f102bc
343c00b3
62d24004
0c56f324
00000804
0336f016
40c3eb96
92c371c3
04c1005c
045c10c3
303c04c9
145c40ac
313c04d1
245c81ac
523c04d9
6006c1ac
853c7c0f
08c30e00
f6bc3fe6
645c09e2
06c30701
0709645c
402c363c
0711045c
81ac303c
0719145c
c1ac313c
08c366f2
09e476bc
39330486
0561245c
245c62c3
323c0569
645c432c
363c0571
045c81ac
103c0579
2007c1ac
145c1c94
21c30201
0209145c
412c313c
0211245c
81ac323c
0219645c
c1ac363c
06356067
045460c7
79dc6107
08c30015
09e476bc
33b30706
642c456c
bbbb601c
bbbb611c
30e406c3
001484dc
0581545c
545c65c3
353c0589
645c432c
363c0591
045c81ac
303c0599
13e4c1ac
c0061394
0565645c
056d645c
0575645c
057d645c
0585645c
058d645c
0595645c
059d645c
050901b3
0565045c
345c6529
a549056d
0575545c
645cc569
045c057d
50c30541
0549045c
42ac303c
0551545c
81ac353c
0559645c
c1ac363c
fff0533c
6f5ca4f7
645c0261
353c0545
64b7420b
02415f5c
054d545c
963cc4d7
9f5c440b
0f5c0227
045c0221
64d70555
64377832
02015f5c
055d545c
7c32686c
100c233c
6d00656c
64cc656f
64cf6d20
aaaa601c
aaaa611c
0006c44f
3c0f042f
1110301c
0000311c
335c6c0c
04c306a4
366417c3
326430c3
62dc6007
145c000c
21c30541
0549145c
412c313c
0551245c
81ac323c
0559545c
c1ac353c
03a1045c
03a9145c
03b1545c
03b9645c
5b946007
402c313c
81ac353c
c1ac963c
01e79f5c
01e10f5c
03c5045c
420b293c
3f5c43b7
345c01c1
693c03cd
c377440b
01a17f5c
03d5745c
183209c3
1f5c0337
145c0181
245c03dd
52c303e1
03e9245c
42ac323c
03f1545c
81ac353c
03f9645c
c1ac363c
5da079c3
613239c3
761423e4
0201045c
045c10c3
303c0209
145c40ac
313c0211
245c81ac
323c0219
60a7c1ac
645c6594
76c30221
0229645c
43ac363c
0231745c
81ac373c
245c04c3
123c0239
d6bcc1ac
0a530a0c
745c5c0c
97c303c1
03c9745c
44ac373c
03d1745c
81ac373c
03d9745c
c1ac373c
6f80e8cc
2f5c6537
245c0281
733c03c5
e2f7420b
01612f5c
03cd245c
733c6517
e2b7440b
01417f5c
03d5745c
58324517
3f5c4277
345c0121
313c03dd
353c402c
763c81ac
e237c1ac
10c30517
1a3517e4
01012f5c
03c5245c
420b573c
6f5ca1f7
645c00e1
073c03cd
01b7440b
00c11f5c
03d5145c
58324217
3f5c4177
345c00a1
08c303dd
09e476bc
09b30006
c00769c3
601c4654
611c11b4
580c0000
14c0353c
3d5423e4
145cebef
21c30781
0789145c
412c313c
0791245c
81ac323c
0799545c
c1ac353c
0010033c
1f5c0137
145c0081
303c0785
60f7420b
00615f5c
078d545c
440b003c
1f5c00b7
145c0041
41170795
40775832
00213f5c
079d345c
00079f5c
0ec0043c
1eb4101c
0014111c
38c324c3
0a5776bc
035c780c
00b30424
76bc08c3
002609e4
c0761596
08040f56
1f36f016
40c3fd96
a2c391c3
20b72006
0bb4301c
0000311c
eebc6c10
30c309f8
60373264
1110301c
0000311c
52892c0c
440c4077
303c0017
082c03c7
5609ac00
341c32c3
6ed20001
0604415c
00013f5c
19c303c3
00213f5c
3ac323c3
70c34664
04c31073
2ac319c3
0a5b5cbc
000770c3
09c37b94
6007600c
30894d54
30a921c3
412c313c
323c50c9
30e981ac
c1ac013c
d528101c
0014111c
089216bc
00070164
40171654
13544007
11544167
10c30017
0d5421c7
618730c3
10c30a54
075421a7
6007744c
4c895154
4e944007
0036c01c
03c36057
03540087
004ac01c
640c19c3
fa80433c
7100502b
002b635c
0383545c
04b465e4
53c37720
301c5364
311c1388
6c0b0000
53e46112
0bc307f4
1abc14c3
e02608e7
801c0533
811c1110
18c30000
6c0c640c
1f3c0c6c
40060080
5abc3ac3
00070a4e
28c3eb94
4097680c
04e4835c
296c04c3
59803cc3
60978664
6097accf
0ccc4d6c
4d8f4800
14c30bc3
08e71abc
19c34097
07c3440f
f8760396
08040f56
0a310abc
00000804
3f36f016
60c3f996
40f7a1c3
1110301c
0000311c
2c106c0c
842c19c3
09f8eebc
326430c3
5a896177
5aa952c3
42ac323c
353cbac9
1ae981ac
c1ac303c
21b72706
03546087
61b76986
353ca157
718003c7
20c30e09
0001241c
11544007
1110301c
0000311c
6eec6c0c
2f5c0ac3
12c300c1
00a14f5c
366424c3
175350c3
14d05ac3
0161065c
065c10c3
303c0169
165c40ac
313c0171
465c81ac
343c0179
72c3c1ac
83e4d2c3
78c30535
d01c83c3
0ac30001
b01c8170
b11c1110
293c0000
40b70180
700c4ac3
146c59c3
31e410c3
60470354
61577994
816743c3
02f32994
59c30026
05f5055c
3fe6748c
03c32037
41172086
2abc6097
2f5c09e0
255c0081
148c05f5
40463f66
09e0bebc
700c4bc3
0bb4501c
0000511c
6f8c540c
2006082c
36644146
326430c3
60076137
0bc3da54
2026600c
00061f5c
2f5c4046
8e6c0025
1cc30006
a19728c3
466435c3
03f250c3
0a13a026
00070dc3
1ac31854
c3c3656c
78a4c884
0161465c
465c04c3
343c0169
065c402c
303c0171
165c81ac
313c0179
73e4c1ac
87c30234
0ac3edf2
0a4066bc
401c09d2
411c0b84
700c0000
2226001c
0bc33664
3a89400c
3aa941c3
422c313c
343c9ac9
8a0c81ac
20c605c3
253cbae9
4664c1ac
06c340c3
40d714c3
0a5e12bc
0dd250c3
66bc04c3
09d20a40
0b84001c
0000011c
001c600c
3664222c
b4dce007
05c3fff6
fc760796
08040f56
3f36f016
40c3e296
b2c361c3
380f2006
a2c34e24
1250d01c
0000d11c
4004923c
f524c9c3
0261145c
145c21c3
313c0269
245c412c
323c0271
145c81ac
313c0279
6af2c1ac
40043a3c
60070486
0023c2dc
0486f324
245c4713
12c301e1
01e9245c
40ac323c
01f1145c
81ac313c
01f9245c
c1ac323c
6d546007
0221145c
145c21c3
313c0229
245c412c
323c0231
145c81ac
313c0239
780fc1ac
67376c2c
03812f5c
0225245c
420b133c
2f5c26f7
245c0361
6717022d
440b133c
1f5c26b7
145c0341
47170235
46775832
03213f5c
023d345c
2df22717
03812f5c
0245245c
345c32c3
12c3024d
0255145c
025d245c
01e1145c
145c21c3
313c01e9
245c412c
323c01f1
145c81ac
313c01f9
133cc1ac
2637fff0
03012f5c
01e5245c
420b113c
2f5c25f7
245c02e1
661701ed
440b133c
1f5c25b7
145c02c1
461701f5
45775832
02a13f5c
01fd345c
200719c3
000c72dc
1893f324
40072bc3
000b82dc
11b4301c
0000311c
67776c0c
b510101c
0014111c
8f6f2f4f
245ccfef
12c302c1
02c9245c
40ac323c
02d1145c
81ac313c
02d9245c
c1ac323c
39546007
678f2757
02c1245c
245c12c3
323c02c9
145c40ac
313c02d1
245c81ac
323c02d9
4facc1ac
47af2757
02c1145c
145c21c3
313c02c9
245c412c
323c02d1
145c81ac
313c02d9
6facc1ac
4f8f4757
02c1145c
145c21c3
313c02c9
245c412c
323c02d1
145c81ac
313c02d9
4757c1ac
03f34faf
03a13f5c
02c5345c
213c2757
4537420b
02812f5c
02cd245c
133c6757
24f7440b
02611f5c
02d5145c
58324757
3f5c44b7
345c0241
275702dd
27af278f
02e1245c
245c12c3
323c02e9
145c40ac
313c02f1
245c81ac
323c02f9
233cc1ac
44770010
02213f5c
02e5345c
420b223c
3f5c4437
345c0201
245702ed
440b213c
2f5c43f7
245c01e1
645702f5
63b77832
01c11f5c
02fd145c
47576186
2026698f
2dc329cf
6c80680c
6757680f
19c36e71
f32422d2
a4bc0757
475709f1
0424025c
20330bd2
40043a3c
60070026
000fc2dc
0026f324
180c1f13
145ca16c
21c301c1
01c9145c
412c313c
01d1245c
81ac323c
01d9145c
c1ac313c
544b63f2
61ec45f2
84dc60c7
61ec000d
6087432c
823c0694
723c00c0
00b30100
0080823c
0180723c
323c540c
3203818c
418c223c
ffff101c
ff00111c
68323183
740f3203
323c542c
3203818c
418c223c
133c3183
1203408c
31c3342f
211c4006
3283ffff
40066077
ffff211c
039432e4
342f1364
e03760cc
23c32226
38bc38c3
540c0a3f
818c323c
223c3203
101c418c
111cffff
3183ff00
32036832
542c740f
818c323c
223c3203
3183418c
32036832
30e3742f
60073364
000812dc
245cf524
12c30141
0149245c
40ac323c
0151145c
81ac313c
0159245c
c1ac323c
0010233c
3f5c4377
345c01a1
223c0145
4337420b
01813f5c
014d345c
213c2357
42f7440b
01612f5c
0155245c
78326357
1f5c62b7
145c0141
5309015d
532912c3
40ac323c
313c3349
536981ac
c1ac323c
fff0233c
3f5c4277
730d0121
420b223c
3f5c4237
732d0101
213c2257
41f7440b
00e12f5c
6257534d
61b77832
00c11f5c
5389336d
53a912c3
40ac323c
313c33c9
53e981ac
c1ac323c
0080233c
2ccc780c
617768a0
00a12f5c
133c538d
2137420b
00812f5c
615753ad
440b133c
1f5c20f7
33cd0061
58324157
3f5c40b7
73ed0041
22d21cc3
180cf324
0a4066bc
580cb733
7f0568cc
580c68cf
6105696c
0006696f
fc761e96
08040f56
0736f016
a1c3fe96
600682c3
12bc6077
30c30a5f
140c5ac3
6b540007
69946007
301c400c
311c1110
8c0c0000
ec6c700c
29e497c3
000ba2dc
72dc4047
503c000b
542bfa80
f889d500
620537c3
21891980
203c61a9
755c00e0
e03704a1
931c97c3
03940004
00534949
445c48a9
113c0564
7f5c41ac
37c30001
30c34664
60073264
000942dc
20178546
408721c3
87c60254
37c3f40b
342b7e05
58896ca0
73c36d20
301c7364
311c1388
6c0b0000
73e46112
301c07f4
311c0bb4
0c0c0000
901c02f3
911c1110
19c30000
6c0c640c
1f3c0c6c
24c30040
5abc38c3
60c30a4e
0bb4801c
0000811c
28c308d2
15c3080c
08e71abc
0b930026
36ec6057
60572c2f
04a4255c
60574def
2cef37ac
57cc6057
60574d0f
0464155c
60572daf
0481255c
01c5235c
155c6057
135c0489
605701cd
0493255c
60574fae
0400033c
0980153c
b0bc4206
605708cb
0500033c
0a80153c
b0bc4206
605708cb
05c4155c
40572f0f
6e20696c
4057696f
61c5696c
29c36b2f
4057680c
04e4335c
296c05c3
366426c3
696c4057
696f6e00
7e204057
605768cf
eccc4d6c
4d8f4b80
040c18c3
1abc15c3
605708e7
680f2ac3
005306c3
02960006
0f56e076
00000804
fb961016
80378086
2fc34077
0a6464bc
08560596
00000804
0136f016
51c340c3
73c362c3
0e00803c
3fe608c3
09e2f6bc
f5244e24
0447353c
135c7180
380f25e4
2604135c
323c3c0f
62d24004
08c3f324
09e476bc
80760006
08040f56
0f36f016
50c3f596
72c361c3
4e24b3c3
005cf524
10c30261
0269055c
40ac303c
0271155c
81ac313c
0279055c
c1ac303c
0400241c
248668f2
22dc4007
f324001c
37d32486
01c33589
313c35a9
15c9402c
81ac303c
a13c35e9
42d2c1ac
7c0cf324
20946087
600778ec
055c1194
10c303c1
03c9055c
40ac303c
03d1155c
81ac313c
03d9255c
c1ac323c
0ac378ef
263c3c2c
363c01c0
54bc0200
24260a07
2c540007
301c31f3
311c106c
6c0c0000
0ac36f0c
253c17c3
366407c0
000710c3
001814dc
03e1055c
055c10c3
303c03e9
155c40ac
313c03f1
255c81ac
323c03f9
0c89c1ac
03c5055c
155c2ca9
4cc903cd
03d5255c
055c0ce9
796c03dd
796f7f05
21c33609
313c3629
5649412c
81ac323c
303c1669
233cc1ac
42b70010
01413f5c
123c760d
2277420b
01212f5c
6297562d
440b033c
0f5c0237
164d0101
38322297
2f5c21f7
566d00e1
10c31689
303c16a9
36c940ac
81ac313c
323c56e9
18ccc1ac
61b76c00
00c11f5c
333c368d
6177420b
00a10f5c
219716ad
440b213c
2f5c4137
56cd0081
78326197
0f5c60f7
16ed0061
39ef3c0c
60877c0c
796c0a94
7b2f7d85
0040973c
833c78ec
07930140
03e1055c
055c10c3
303c03e9
155c40ac
313c03f1
255c81ac
323c03f9
6c49c1ac
60872a06
000f94dc
7b05796c
973c7b2f
155c0040
21c303e1
03e9155c
412c313c
03f1255c
81ac323c
03f9055c
c1ac303c
0080833c
155c7b0f
21c303c1
03c9155c
412c313c
03d1255c
81ac323c
03d9055c
c1ac303c
78cc78ef
78cf6105
3509996c
352921c3
412c313c
85ac233c
78cc500f
800c133c
818c323c
223c3203
001c418c
011cffff
3083ff00
32036832
313c700f
3103818c
418c213c
68323083
702f3203
01c1255c
255c02c3
323c01c9
055c402c
303c01d1
155c81ac
313c01d9
64d2c1ac
60c77c0c
78cc2a94
00079f5c
222606c3
38c323c3
0a3f38bc
13c330e3
25f21364
ffff101c
0000111c
323c502c
3203818c
418c223c
ffff001c
ff00011c
68323083
21c33203
323c23a3
3203818c
418c223c
68323083
702f3203
0e00ba3c
3fe60bc3
09e2f6bc
60877c0c
5c2c3b94
0161055c
055c10c3
303c0169
155c40ac
313c0171
055c81ac
403c0179
155cc1ac
01c30181
0189155c
402c313c
0191055c
81ac303c
0199155c
c1ac313c
60066037
0011311c
055c6077
10c301a1
01a9055c
40ac303c
01b1155c
81ac313c
01b9055c
c1ac303c
0ac360b7
34c316c3
0a22a0bc
18c30533
3a8f240c
482c28c3
38c35aaf
7acf6c4c
006c08c3
19c31aef
3a0f240c
482c29c3
39c35a2f
7a4f6c4c
006c09c3
301c1a6f
311c106c
6c0c0000
1ac3b8cc
31a4115c
8e4c2037
16c30ac3
35c34226
0bc34664
09e476bc
01c32006
f0760b96
08040f56
0336f016
80c3fe96
72c351c3
440c93c3
1110301c
0000311c
640c2c0c
40c30c6c
035424e4
31944047
c5867c0c
02546087
756cc806
802654cc
00064f5c
0f5c0046
866c0025
13c30006
466436c3
06f240c3
66bc05c3
00260a40
05c30593
0a4066bc
301c09d2
311c0b84
6c0c0000
2228001c
301c3664
311c1110
6c0c0000
04c36e0c
5c0c2226
50c33664
15c308c3
39c327c3
0a6280bc
05c30dd2
0a4066bc
301c09d2
311c0b84
6c0c0000
222d001c
00063664
c0760296
08040f56
fd961016
305c40c3
60071ce4
301c1d94
311c1100
6c0c0000
0090233c
141d6146
402c3230
60776037
60b76026
03a0021c
201c12c3
211cc9cc
34c30014
09f3c8bc
345c6026
03961ce7
08040856
01fc021c
0100101c
bebc4006
080409e0
f7967016
1b64505c
1b44405c
800734c3
000d02dc
0a01045c
045c10c3
303c0a09
145c40ac
313c0a11
245c81ac
323c0a19
17f3c1ac
d2dc6007
045c0009
10c30201
0209045c
40ac303c
0211145c
81ac313c
0219245c
c1ac323c
b4dc60a7
145c0008
21c306c1
06c9145c
412c313c
06d1245c
81ac323c
06d9045c
c1ac303c
79546007
fff0233c
3f5c41f7
345c00e1
123c06c5
21b7420b
00c12f5c
06cd245c
033c61d7
0177440b
00a10f5c
06d5045c
383221d7
2f5c2137
245c0081
61d706dd
59946007
06e1045c
045c10c3
303c06e9
145c40ac
313c06f1
245c81ac
323c06f9
133cc1ac
22370010
01012f5c
06e5245c
420b013c
1f5c00f7
145c0061
421706ed
440b323c
3f5c60b7
345c0041
021706f5
00771832
00211f5c
06fd145c
4c0c780c
02176909
13e410c3
48e92334
2f5c4037
245c0001
600606c5
06cd345c
06d5345c
06dd345c
0221045c
045c10c3
303c0229
145c40ac
313c0231
245c81ac
323c0239
04c3c1ac
fff0133c
0a0cd6bc
04c30093
0a1316bc
0861045c
045c10c3
303c0869
145c40ac
313c0871
245c81ac
423c0879
045cc1ac
10c30a01
0a09045c
40ac303c
0a11145c
81ac313c
0a19245c
c1ac323c
00b3bfe5
106c601c
0000611c
d4dca007
0996fff3
08040e56
3f36f016
c0c3f496
256c41c3
921c91c3
09c30004
323c400c
3203818c
418c223c
ffff501c
ff00511c
68323583
600f3203
263c61c3
86c3044e
818c323c
223c3203
3583418c
32036832
71c3780f
064e273c
818c323c
223c3203
3583418c
32036832
61c37c0f
084e263c
818c323c
223c3203
3583418c
32036832
31c3780f
0a4e233c
323ca3c3
3203818c
418c223c
68323583
0ac33203
51c3600f
0c4e253c
818c323c
223c3203
101c418c
111cffff
3183ff00
32036832
29c3740f
40f7480b
7fe532c3
51b46027
280c28c3
808c013c
5c0c00b7
808c323c
81acd13c
b23c382b
70ec80ac
3c3c64f2
70ef4a80
40774e24
3cc3f524
23a4135c
203724f2
011321c3
005c0cc3
003723c4
235c3cc3
005723e4
341c30c3
60770400
f32462d2
19542007
0077140c
0854b2e4
00070bc3
60571294
02e403c3
50ec0e94
60974077
686c03c3
059403e4
30c3088c
0354d3e4
16640017
4cac70ec
0d94b2e4
315c1cc3
65d22384
14c30cc3
20933664
66bc04c3
20130a40
03c360d7
24dc0027
740c0008
7e9432e4
680c29c3
011c0006
3083ffff
680f6172
686c50ec
333c292b
28c380ac
50ec680f
096b688c
802c333c
70ec7c0f
20976cac
80ac333c
2ac3780f
7411a811
4c0c39c3
818c323c
223c3203
001c418c
011cffff
3083ff00
32036832
640f19c3
4c0c38c3
818c323c
223c3203
3083418c
32036832
640f18c3
323c5c0c
3203818c
418c223c
68323083
7c0f3203
323c580c
3203818c
418c223c
68323083
780f3203
4c0c3ac3
818c323c
223c3203
3083418c
32036832
600f0ac3
323c540c
3203818c
418c223c
ffff101c
ff00111c
68323183
740f3203
50cf4386
6d00716c
cf5c718f
60c60147
82376137
a1b7a097
00e7df5c
62f770ec
0f3c6e0c
36640100
04c30093
0a4066bc
408c3b3c
033c3b84
303c01f4
6cc30f30
3a1d163c
045321c3
3be4690c
c0971c94
a951c92f
106c301c
0000311c
6c0c6c0c
682f6c29
084f0006
296f30ec
f5246e24
03d2098c
a98fa006
0400341c
3c546007
0753f324
21e448ac
40073c54
0733de94
303c0cc3
4ccc5a1d
60976911
a951692f
106c301c
0000311c
6c0c6c0c
682f6c29
b0ec284f
01c3a96f
802c03f3
c02fc006
21b72097
00e7df5c
0147cf5c
0237c137
42f740ec
c92c60cc
31e416c3
2cc30835
1284325c
e8bc65f2
00930a0a
05c36a0c
04c33664
5f3c0073
00070100
0213df94
0f30503c
100c353c
265c6cc3
0cc32304
26643980
000610c3
ee942007
0c96f753
0f56fc76
00000804
0736f016
50c3fc96
13e4705c
0000801c
a01c48c3
a11c106c
9f3c0000
12b300c0
60077c0c
0008f2dc
100c683c
1444355c
680c4f00
62dc6007
83d20008
03356027
680f7fe5
1444355c
60076f01
80077b94
055c7994
19c306e4
34c34486
0a4e5abc
70940007
410660d7
40d74ccf
6105696c
40d7698f
1404355c
28ef2f01
8d6c60d7
0684355c
0a946027
111c2006
300f1200
502f5c0c
0687355c
60060153
1600311c
3c0c700f
4046302f
0687255c
103c100c
502c808c
341c30c3
2c80ffff
808c323c
241c6580
6d00ffff
808c233c
ffff341c
233c6d00
341c808c
6d00ffff
341c33e3
30a3ffff
60d7700f
2def2086
5c0c60d7
500c4d0f
818c323c
223c3203
101c418c
111cffff
3183ff00
32036832
502c700f
818c323c
223c3203
3183418c
32036832
7c0c702f
40374026
111c2006
20770002
40b74006
20d705c3
600623c3
0a22a0bc
e0858026
0001821c
640c1ac3
6de96c0c
70dc83e4
0496fff6
0f56e076
00000804
01fc021c
40062026
09e0bebc
00000804
0336f016
505c60c3
e0062284
833c6e24
901c4004
911c106c
0e330000
6007742c
7fe56c54
6007742f
752c6894
754c6af2
544c68f2
600c09c3
6d296c0c
509423e4
54ecf524
17544007
51e434ac
00060494
0153080f
35e4680c
280f0294
34cc54ac
74cc28cf
365c4caf
7fe522a4
22a7365c
54ef4006
52e4546c
00060594
2287065c
348c0193
748c288f
365c4c6f
35e42284
746c0494
2287365c
2284365c
746f6ed2
2284365c
148f0c8c
2284365c
ac6f6c8c
2284365c
00b3ac8f
2287565c
b48fb46f
2006158c
28c3358f
f32449d2
802c00f3
602f6006
0a0ae8bc
1af204c3
323c01d3
744f0010
600c09c3
6d496c0c
06c3742f
556c350c
0a68c8bc
e025b46c
22a4165c
72e421c3
c0768c14
08040f56
0f36f016
b0c3f796
92c3a1c3
06e4005c
02001f3c
60064206
0a4e5abc
000780c3
0009e4dc
2cf16217
23866217
42172ccf
6c80696c
6217698f
201c2d6c
211c0800
440f0001
602641c3
0604311c
027e343c
621701c3
686c4cec
333ca92b
303c82ac
51c3047e
4cec6217
c96b688c
832c333c
067e353c
621761c3
6cac6cec
363c7012
71c3087e
0a7e873c
a23c21c3
82c30c7e
323c440c
3203818c
418ca23c
ffff201c
ff00211c
68323283
640f3a03
323c500c
3203818c
418c223c
ffff101c
ff00111c
68323183
700f3203
323c400c
3203818c
418c223c
68323183
600f3203
323c540c
3203818c
418c223c
68323183
740f3203
323c580c
3203818c
418c223c
68323183
780f3203
323c5c0c
3203818c
418c223c
68323183
7c0f3203
440c18c3
818c323c
223c3203
501c418c
511cffff
3583ff00
32036832
bf5c640f
c0a600c7
2217c037
201c2137
211cffff
40b70000
60f77fe6
00e79f5c
760c59c3
36640fc3
f0760996
08040f56
0336f016
70c3fe96
1074001c
0000011c
f6bc3fe6
c00609e2
10a8801c
0000811c
106c901c
0000911c
640c18c3
06e92f00
32540007
035400a7
2e940027
6c4c650c
2a9437e4
600764ec
66c92594
07c365f2
0a096cbc
39c30433
a58c4c0c
0056303c
7f327fe5
8b2c6037
402607c3
466435c3
640c18c3
4ec96f00
3fe512c3
2f5c2077
4ecd0021
640c18c3
275c6f00
4cef3164
7fe50073
c68564ef
0340631c
001cc694
011c1074
76bc0000
029609e4
0f56c076
00000804
50c3f016
1074001c
0000011c
f6bc3fe6
000609e2
10a8401c
0000411c
106c601c
0000611c
4c00700c
20072ae9
6b692954
26946007
6c4c690c
229435e4
08942047
64f268ec
eaede066
7fe50373
20870313
28ec1294
fff0313c
11942007
eaede0a6
6c00700c
700c2cef
780c4c00
2e896c0c
00d32acd
04942067
602568ec
068568ef
0340031c
001cd094
011c1074
76bc0000
0f5609e4
00000804
50c33016
f5246e24
1c04105c
205c4006
205c1c07
205c1c27
341c1c47
6ad20400
0113f324
6006842c
05c3642f
0a269ebc
39f214c3
08040c56
40c33016
533c6e24
01b34004
642cf524
22c7345c
345c63f2
a2d222e7
04c3f324
0a65d0bc
22c4145c
0c5632f2
00000804
ffffffff
ffffffff
ffffffff
feffffff
ffffffff
ffffffff
ffffffff
ffffffff
ffffffff
ffffffff
00000000
00000000
01000000
ffffffff
01000000
00000000
00000000
00000000
ffffffff
ffffffff
ffffffff
00000001
00000000
00000000
00000000
00000000
00000000
00000000
00000000
204c5353
656d6974
00000072
4641544f
50435420
636f5320
0074656b
0336f016
1114301c
0000311c
ac0c6c0c
0b08301c
0000311c
60076c2c
301c5a94
311c0b84
6c0c0000
2119001c
0a333664
640c19c3
100462f2
29c37fe5
702c680f
62f2682f
f02b684f
cca9740c
1194c007
640c18c3
0404335c
14c305c3
1fe73664
740c0854
05c7203c
68802c0c
02d6635c
341c7381
331cf000
23945000
200675ac
0008111c
60073183
28c31654
335c680c
05c30424
366414c3
1fe720c3
18c30954
335c640c
05c30444
366414c3
28c30353
0073680c
640c18c3
04c36dcc
02333664
680c28c3
0484335c
14c305c3
01333664
0b08901c
0000911c
1114801c
0000811c
8c2c39c3
a5948007
0bb4301c
0000311c
00266c0c
1341135c
0872b8bc
0f56c076
00000804
ff96f016
301c50c3
311c1114
2c0c0000
040cc46c
6109400c
68d26037
942b744c
6de96e00
62d26037
68a9402c
13546027
11546067
15c385ac
00017f5c
466437c3
301c0af2
311c0bb4
0c0c0000
1abc15c3
051308e7
742f6006
f5248e24
78bc0046
788c08cc
78ac64d2
0053ac2f
b8afb88f
1114301c
0000311c
4c6c6c0c
6025686c
0046686f
08cc82bc
4004343c
f32462d2
20660046
0fe4301c
0000311c
d4bc4d0c
019608c8
08040f56
0f36f016
201cff96
211c1114
680c0000
cc6cec0c
933c6e24
82c34004
0ef0b01c
0000b11c
0bb4a01c
0000a11c
0026f524
08cc78bc
69f2780c
82bc0026
09c308cc
49540007
08f3f324
340cb82c
7fe5382f
0026780f
08cc82bc
42d229c3
355cf324
608701d1
08c30994
335c600c
07c304e4
366415c3
548cfb93
31c32889
89806205
6c0c7c0c
0010033c
0060143c
eabc40c6
38c308cb
303c4c0c
33c40b0d
f88c133c
696c2037
14c307c3
00014f5c
366424c3
5fe720c3
18c30854
6d8c640c
15c307c3
f6b33664
680c2bc3
100c4ac3
0040153c
f5b33664
0bb4301c
0000311c
02e66c0c
1341135c
0872b8bc
f0760196
08040f56
301c1016
311c0bb4
8c0c0000
6d0c71cc
200604c3
02e63664
1341145c
0872a2bc
08040856
126410c3
ff32001c
31b42067
0608201c
4130211c
680c680c
0400341c
ff34001c
25946007
680c28f2
680f6a72
341c680c
03330400
08942027
6b72680c
680c680f
0800341c
20470213
680c0894
680f6c72
341c680c
00f31000
6d72680c
680c680f
2000341c
63f20006
ff35001c
00000804
0608301c
4130311c
341c6c0c
60070400
201c1194
211c0620
680c2040
0054033c
301c1df2
311c0620
6c0c2040
0001341c
001c63f2
0804ff35
40c31016
0a6c34bc
0608301c
4130311c
341c6c0c
001c0800
6007ff2f
301c4394
311c0628
6c0c2040
0001341c
ff34001c
38546007
0600301c
2040311c
4c0f4046
0620101c
2040111c
341c640c
60070001
640c2754
0004341c
22946007
01c323c3
600c2505
0080341c
640c7dd2
40857161
04a8231c
201cf794
211c0620
680c2040
0002341c
301c7dd2
311c0620
6c0c2040
0002341c
ff35001c
000665d2
001c0073
0856ff33
00000804
40c31016
0a6c34bc
0628301c
2040311c
341c6c0c
001c0002
6007ff34
301c4054
311c0600
40862040
101c4c0f
111c0620
640c2040
0001341c
2d546007
3283640c
29946007
01c323c3
600c2485
0040341c
71017dd2
4085640f
04a8231c
201cf794
211c0620
680c2040
0002341c
680c65f2
0004341c
201c79d2
211c0620
680c2040
0005341c
680c6bd2
0004341c
ff31001c
00b365d2
ff33001c
00060053
08040856
50c37016
41c363c3
12c34264
301c1364
311c0608
6c0c4130
1000341c
ff2f001c
66946007
0100131c
001c0654
131cff32
5e940080
0628301c
2040311c
341c6c0c
001c0004
6007ff34
301c5354
311c060c
40262040
301c4c0f
311c0604
8c0f2040
308c213c
4c0f6085
0600301c
2040311c
4c0f4206
0620201c
2040211c
341c680c
60070001
680c3354
0004341c
2e946007
288c013c
42c313c3
01334405
341c700c
7dd20010
1a1d353c
2025680f
f71410e4
001c4006
011c0620
101c2040
111c0648
600c2040
0080341c
640c7dd2
40857961
f8944587
0620201c
2040211c
341c680c
60470003
0006fc94
001c0073
0e56ff33
00000804
0620201c
2040211c
341c680c
7dd20002
0408201c
2040211c
0408101c
2040111c
341c680c
79f20004
60876069
63660994
301c640f
311c0500
40662040
61460113
301c640f
311c0500
40262040
201c4c0f
211c0520
680c2040
0008341c
00067dd2
00000804
ff96f016
71c360c3
226413c3
301c4037
311c0628
6c0c2040
0008341c
ff34001c
52dc6007
3f5c0011
30640001
34e48006
60170815
241c23c3
4037007f
0100401c
60877869
a0860954
07546047
640f6006
ff32001c
a1061f93
100c353c
4017640f
602732c3
301c1394
311c0608
6c0c4130
2000341c
ff2f001c
94dc6007
301c000e
311c060c
40172040
601702f3
16946007
0794a107
0408301c
2040311c
4c0f4026
060c301c
2040311c
4c0f4006
0500301c
2040311c
4c0f4026
001c04d3
6017ff30
404723c3
000c44dc
060c301c
2040311c
4c0f4006
0c94a107
0155343c
0408201c
2040211c
0004680f
01d5343c
34c30173
201c6272
211c0408
680f2040
343c0004
680f00c5
0600301c
2040311c
4c0f4806
0620101c
2040111c
341c640c
60070001
000922dc
341c640c
60070004
0008c4dc
01c323c3
600c2485
0040341c
79017dd2
4085640f
f8944587
32c34017
1e946027
400617c3
0620401c
2040411c
0664001c
2040011c
341c700c
7dd20020
313c600c
4025027f
f71425e4
0620201c
2040211c
341c680c
7dd20002
40170c33
23944007
00871869
301c0794
311c0500
40662040
00470113
301c0794
311c0500
40262040
201c4c0f
211c0620
680c2040
0002341c
201c7dd2
211c0520
680c2040
0008341c
07937dd2
ff35001c
23c36017
37944047
0620201c
2040211c
341c680c
7dd20002
0408201c
2040211c
0408101c
2040111c
341c680c
79f20004
60877869
343c0a94
640f01b5
0500301c
2040311c
01334066
00a5343c
301c640f
311c0500
40262040
201c4c0f
211c0520
680c2040
0008341c
00937dd2
ff33001c
00060053
0f560196
00000804
0f36f016
12c3a1c3
c25783c3
526450c3
0024353c
62f24406
723c4206
973c108c
141d100c
423cb690
341d180c
001c2620
4007ff32
000b84dc
0044353c
2e546007
0100431c
301c0c94
311c0408
40262040
321c4c0f
201c00f8
01530083
0408301c
2040311c
321c4c0f
201c00f8
4c0f0081
400648c3
0520601c
2040611c
0540001c
2040011c
341c780c
64070028
343cfc94
600f024f
27e44025
301cf614
311c0508
40062040
301c4c0f
311c0504
40462040
201c4c0f
211c0520
680c2040
0001341c
301c7df2
311c0508
40262040
201c4c0f
211c0520
680c2040
0040341c
640c7dd2
0544201c
2040211c
642c680f
644c680f
646c680f
353c680f
201c0084
211c0520
60072040
1ac31094
501c8006
511c0520
801c2040
811c0544
601c2040
611c0548
07d32040
341c680c
7dd20040
201c648c
211c0544
680f2040
680f64ac
680f64cc
680f64ec
343cfc33
65f20034
341c740c
ff930040
400601c3
0034323c
740c65f2
0040341c
a03cff93
38c3024f
40254c11
f31427e4
20c30006
0034303c
740c66f2
0080341c
40067dd2
62975810
2b9da33c
07e40025
40250334
8025fe13
4be41984
0006d314
0f56f076
00000804
3f36f016
81c3fb96
43c3b2c3
cf5cc457
50c30284
1cc35264
0f3c27d2
24d70080
b0bc4186
353c08cb
44060024
420662f2
108ca23c
100c9a3c
7690141d
123ce037
341d180c
001c2620
4007ff32
000e54dc
0044353c
2f546007
0100131c
301c0d94
311c0408
e0262040
321cec0f
101c00f8
2c0f0083
301c0173
311c0408
4c0f2040
00f8321c
0081201c
24174c0f
601c4006
611c0520
001c2040
011c0540
780c2040
0028341c
fc946407
024f313c
4025600f
f6142ae4
0508301c
2040311c
ec0fe006
0014153c
301c28d2
311c0504
40462040
00f34c0f
0504301c
2040311c
ec0fe026
0520201c
2040211c
341c680c
7df20001
0104353c
301c68d2
311c0508
40262040
00f34c0f
0508301c
2040311c
ec0fe046
1c542007
0520201c
2040211c
341c680c
7dd20040
201c700c
211c0544
680f2040
680f702c
680f704c
680f706c
0084353c
0520201c
2040211c
e4976af2
801c68c3
d01c0000
d11c0548
0b332040
341c680c
7dd20040
201c708c
211c0544
680f2040
680f70ac
680f70cc
680f70ec
1cc3fcf3
bf5c23d2
06c30027
323c4006
69f20034
0520101c
2040111c
341c640c
ff130040
66d23cc3
00401f3c
2a1d313c
600c0053
0544101c
2040111c
4025640f
2ae40085
56c3e514
17c347c3
303c0006
69f20034
0520201c
2040211c
341c680c
ff130080
67d23cc3
4c0c3dc3
3203740c
0093700f
680c2dc3
0025640f
8085a085
0ae42085
821ce514
79840001
b9846984
21c32017
b61482e4
05960006
0f56fc76
00000804
60061016
413c00d3
403c3a1d
60253b9d
fa1432e4
08040856
60061016
413c00d3
403c359d
6025371d
fa1432e4
08040856
0136f016
71c380c3
63c342c3
43e70006
640615b4
0006ad20
01d310c3
1a1d273c
400d323c
38c303a3
1b9d033c
508d023c
04c382f2
16e42025
8076f214
08040f56
60c37016
136441c3
036402c3
128d303c
5032780f
128d523c
808c343c
028d133c
223c06c3
203c328d
b480027e
063451e4
111c2006
68800001
253c600f
380c800c
780f6880
043432e4
6025600c
353c600f
400c808c
600f6d00
08040e56
32c33016
62125fe5
01807f85
01d32580
640c800c
033543e4
01730026
3f851f85
033443e4
00b31fe6
40075fe5
0006f215
08040c56
1f36f016
80c3fe96
72c3a1c3
cf5c93c3
42c30184
24544007
64c38006
03d354c3
17c30fc3
4e8139c3
0a70e8bc
66811ac3
38c34e20
34e34ee1
23e40006
00260235
68a02017
6ae128c3
22e34017
023532e4
40570025
c0258100
6ce4a085
04c3e214
f8760296
08040f56
0f36f016
91c3a0c3
73c382c3
60c30006
029340c3
660119c3
30e3ac20
460118c3
53e412e3
352007b4
002632e3
02b413e4
3ac30006
c0252e61
67e48085
f076ec14
08040f56
50c3f016
23c342c3
83e70006
64061ab4
623cee20
323cfff0
7f85100c
55802580
01b30006
353ca40c
03a3408d
04c3080f
053c83d2
dfe5700d
5f853f85
f315c007
08040f56
0f36f016
92c3b0c3
808c023c
442c840c
808c623c
ffff101c
0000111c
03e431c3
303c0754
141d0010
63c33230
79c36364
163c7364
313c728d
91a0800c
43e433e3
5fe50235
808c313c
363c49a0
29a0028d
800c273c
82c4a2e3
0173b120
02355ae4
24203fe5
0010363c
636463c3
48845884
f5b410e4
039410e4
f13442e4
536451c3
ffff201c
0000211c
03e432c3
243c0c54
313c808c
4980800c
0010303c
3230141d
536453c3
728d353c
028d053c
33e351a0
023523e4
303c3fe5
49a0800c
23e433e3
3fe50235
808c303c
49e325a0
29a40133
023524e4
353c3fe5
53c30010
38f25364
f63429e4
800c363c
4bc37580
f076700f
08040f56
00b36006
203c4006
60253b9d
fb1431e4
00000804
000630c3
002566d2
03540407
ff736132
00000804
213c31c3
6212fff0
01807f85
303c00b3
64f2fe4f
40075fe5
023cfb15
08040010
3f36f016
c0c3fa96
b2c320b7
9f5c83c3
09c30224
36bc2497
70c30a72
02dc0007
303c000b
a33c100c
29c3ffc0
09813ac3
0a722cbc
d3c36406
501cd0a4
511c13a0
140c0000
22bc17c3
940c0a72
1bc304c3
38c32dc3
0a70c8bc
043c38c3
401c3b9d
411c13a4
100c0000
2dc319c3
c8bc37c3
700c0a70
6d012ac3
0cc360f7
22bc18c3
98c30a72
893c97a4
c884100c
0087cf5c
6b8029c3
100c633c
602537c4
b33c39a4
c5c3130c
23c360d7
40774025
60d70b13
5fe723c3
2cc30694
4f01680c
01534177
680c2cc3
01400f3c
2d002bc3
a8bc4057
2cc30a71
af00680c
38845410
13a4201c
0000211c
e037880c
13c303c3
34c34157
0a7130bc
68202ac3
02b3740f
60256157
2cc36177
8f00680c
3884b00c
13c303c3
13a4301c
0000311c
37c34c0c
0a7164bc
700f7420
080c2cc3
60076301
0884e894
13a4301c
0000311c
27c32c0c
0a7116bc
dd150007
41576117
fe7f233c
921c6137
821cffff
df85fffc
fffcb21c
0000931c
0097a715
22bc2497
00970a72
13a0301c
0000311c
2dc32c0c
86bc37c3
06960a71
0f56fc76
00000804
0736f016
70c3fe96
92c381c3
a01c63c3
a11c10f8
2ac30000
8c0c680c
0400001c
21c32006
27cc301c
0015311c
50c34664
14540007
6297c037
17c36077
39c328c3
0a7246bc
680c2ac3
05c38c4c
21c32006
27cc301c
0015311c
02964664
0f56e076
00000804
60c37016
42c351c3
22bc12c3
343c0a72
53e4280c
153c0934
253c288c
602601f4
363c3223
0e561b9d
00000804
ff961016
f88c213c
41524880
60062080
81a20133
84098037
4f5c81a1
840d0001
3fe56025
f67432e4
08560196
00000804
25001016
00936006
81a18409
3fe56025
fb7432e4
08040856
031cff96
17b40200
0200231c
131c14b4
11b40200
0076303c
0b0d333c
fff0233c
0076313c
0b0d333c
32a37fe5
f88c233c
00734037
60376026
00011f5c
019601c3
00000804
201c6026
211c0404
680e4101
13a8201c
0000211c
0804680d
3f36f016
60c3fb96
92c320b7
0f5cc3c3
00770261
13a0301c
0000311c
2c0f2006
13a4301c
0000311c
60062c0f
4140311c
4000201c
c31c4c0f
08b40100
0001b01c
10c30097
0100131c
b01c0335
3b3c0002
60250817
100c533c
10f8801c
0000811c
680c28c3
05c38c0c
21c32006
27c0301c
0015311c
00f74664
608608f2
4140311c
4000001c
04330c0f
9cbc15c3
3b3c08cb
60250857
100c733c
640c18c3
07c38c0c
21c32006
27c0301c
0015311c
301c4664
311c13a0
0c0f0000
11940007
311c6086
201c4140
4c0f4000
0b84301c
0000311c
001c6c0c
36642221
30b30026
9cbc17c3
08c308cb
8c0c600c
200607c3
301c21c3
311c27c0
46640015
13a4801c
0000811c
040f18c3
db540007
9cbc17c3
06c308cb
52bc2097
09c30a73
52bc1cc3
db3c0a73
06c3300c
36bc1dc3
40c30a72
100c303c
19817f85
0a722cbc
fe00203c
280c343c
a384a2c3
00105d3c
040c18c3
2a3c19c3
35c301f4
0a70c8bc
288c3a3c
2c3c6212
20d70030
38c30580
42322c0c
0a70b0bc
040c18c3
9cbc17c3
09c308cb
100c153c
08cb9cbc
380c7b3c
09c38037
27c320d7
0abc36c3
001c0a73
011c0a00
16c34101
bcbc27c3
001c0a70
011c0200
19c34101
bcbc27c3
001c0a70
011c0800
19c34101
bcbc27c3
06c30a70
12c34097
9cbc2085
645708cb
12946007
9abc0417
3f3c0bae
033c0140
0417fe7e
23c316c3
0bae9ebc
211706c3
0a7352bc
06c300d3
44572417
0a736abc
400c3b3c
fff0233c
035c7980
05f2fff9
7fe55fe5
fa154007
0400101c
4101111c
440e4006
fff02a3c
7fff231c
640b0535
30a31f06
640b00b3
323c3364
336419ac
323c640e
501c0acb
511c0406
740e4101
0400201c
4101211c
3364680b
680e6272
1dc306c3
0a7236bc
303c40c3
7f85100c
2cbc1981
203c0a72
343cfe00
0980280c
0402101c
4101111c
440e40a6
3364640b
ffe0203c
19ac323c
640e3364
13c3740b
303c1364
341cfff0
40460800
23c362f2
401c21a3
411c0406
500e4101
0600001c
4101011c
27c316c3
0a70bcbc
3364700b
700e6272
60076057
201c1854
211c0402
680b4101
6e723364
680b680e
61723364
301c680e
311c13a8
00060000
23c30c0d
68091404
01d37ed2
0402301c
4101311c
23644c0b
4c0e4172
680b23c3
60073164
301cfd15
311c0402
40064101
201c4c0e
211c0202
60064101
016f323c
0400001c
4101011c
21e410c3
301cf794
311c0200
00264101
680b0c0e
fffc341c
680e6072
341c680b
7dd24000
20970497
08cb9cbc
20060497
4101111c
6abc4097
401c0a73
411c10f8
700c0000
00d7ac4c
21c32006
27c0301c
0015311c
700c5664
301cac4c
311c13a0
0c0c0000
21c32006
27c0301c
0015311c
700c5664
301c8c4c
311c13a4
0c0c0000
21c32006
27c0301c
0015311c
60864664
4140311c
4000101c
00062c0f
fc760596
08040f56
1f36f016
b0c3f896
a2c391c3
9abcc3c3
01f70bae
9abc0ac3
01b70bae
9abc09c3
20c30bae
10f8301c
0000311c
6eec6c0c
219701d7
30c33664
60073264
000c94dc
41d76197
0200331c
000c35dc
0200231c
000bf5dc
0100331c
501c06b4
231c0104
03350100
0204501c
22dc60e7
40e7000b
000af2dc
10f8801c
0000811c
680c28c3
05c38c0c
21c32006
2798301c
0015311c
60c34664
1a540007
600c08c3
05c38c0c
21c32006
2798301c
0015311c
70c34664
15940007
640c18c3
06c38c4c
27c317c3
2798301c
0015311c
301c4664
311c0b84
6c0c0000
2221001c
0f533664
15c306c3
08cb9cbc
15c307c3
08cb9cbc
17c30bc3
01c02f3c
0bae9ebc
16c30ac3
01802f3c
0bae9ebc
131c2197
05b40100
531ca1d7
1c350100
10f8301c
0000311c
9f5c4c0c
00060007
c0b70077
10fc301c
0000311c
0c896c0c
00650f5c
06c38aac
61d727c3
01374664
00811f5c
38c30313
9f5c4c0c
00060007
c0b70077
10fc301c
0000311c
0c896c0c
00650f5c
06c38a8c
35c327c3
01774664
00a11f5c
826481c3
16c30cc3
92bc4197
00070bae
301c0915
311c0b84
6c0c0000
2204001c
501c3664
511c10f8
740c0000
06c38c4c
21c32006
2798301c
0015311c
740c4664
07c38c4c
21c32006
2798301c
0015311c
08c34664
00260053
f8760896
08040f56
3f36f016
01b7f696
417791c3
af5c83c3
df5c02c4
301c02e4
311c10f8
6c0c0000
01c36eec
28c31ac3
30c33664
62773264
60070026
000b54dc
01210f5c
931c30c3
02350100
40066026
0100831c
40260235
02a303c3
1f5c0137
c1c30081
2cc3c264
501c46f2
a31c0104
03350100
0204501c
10f8b01c
0000b11c
600c0bc3
05c38c0c
21c32006
27ac301c
0015311c
70c34664
1bc30ed2
8c0c640c
200605c3
301c21c3
311c27ac
46640015
0bf260c3
0b84301c
0000311c
001c6c0c
36642221
0e130026
101c0dc3
9cbc00c0
07c308cb
9cbc15c3
06c308cb
9cbc15c3
07c308cb
2ac32557
08cbb0bc
219706c3
b0bc29c3
2cc308cb
a31c44f2
1e350100
10f8301c
0000311c
01574c0c
8f5c0037
df5c0027
301c0047
311c10fc
6c0c0000
1f5c2c89
8aac0065
1ac307c3
39c326c3
01f74664
00e12f5c
3bc30353
01574c0c
8f5c0037
df5c0027
301c0047
311c10fc
6c0c0000
1f5c2c89
8a8c0065
1ac307c3
39c326c3
02374664
01012f5c
826482c3
10f8501c
0000511c
8c4c740c
200607c3
301c21c3
311c27ac
46640015
8c4c740c
200606c3
301c21c3
311c27ac
46640015
4c116617
0a9608c3
0f56fc76
00000804
333c30c3
333c080d
03c30b8d
00000804
40c31016
34c34364
ff00341c
301c6bd2
311c0b84
6c0c0000
222f001c
441c3664
301c00ff
311c0b84
6c0c0000
051c04c3
36648200
08040856
ff961016
000620c3
303c00b3
201700a7
323c0580
133c009f
2037fd00
00013f5c
f4356127
08560196
00000804
ff963016
400640c3
013302c3
00a7303c
0c807a05
0010323c
236423c3
513c3122
a037fd00
00013f5c
f1356127
0c560196
00000804
fe967016
326430c3
12646077
0bb4301c
0000311c
2027cc0c
28d21954
28542047
20678006
000a24dc
182c0693
40bc4026
40c308e6
80074264
301c3c94
311c0b84
6c0c0000
2122001c
182c0233
40662006
08e640bc
426440c3
2b948007
0b84301c
0000311c
001c6c0c
36642123
182c0fd3
41062006
08e640bc
426440c3
19948007
0b84301c
0000311c
001c6c0c
fdd32124
2006182c
40bc4186
40c308e6
89f24264
0b84301c
0000311c
001c6c0c
fbd32125
0bb4201c
0000211c
ae0c682c
6ccc786c
200602c3
40c33664
4f540007
0110101c
08cb9cbc
1000143c
6057308f
408723c3
3f5c3394
345c0021
640c01d5
323c4057
640f231b
1110301c
0000311c
6c0c6c0c
60276f0b
355c0554
60270c99
60260594
516664cd
60260093
400664cd
355c450d
60070a89
255c2254
32c30301
0309255c
41ac323c
60276037
3f5c1894
64cd0001
450d5166
60570253
2f5c68f2
245c0021
640c01d5
00d34057
345c60a6
640c01d5
323c40a6
640f231b
029604c3
08040e56
1f36f016
83c3ff96
0164cf5c
636460c3
536452c3
0181af5c
0bb4301c
0000311c
2ac36c10
93c36500
2bc39364
9f5c686c
8fcc0007
16c30bc3
35c34006
70c34664
301c0af2
311c0b84
6c0c0000
211f001c
14133664
315c1bc3
606517c4
32835f86
c3878180
631c0b54
08540089
0654c287
0454c827
00a1631c
301c0a94
311c1118
6c0c0000
06c36dec
366414c3
00e6631c
631c0d54
0a5400e2
00db631c
631c0754
045400e4
00e7631c
18c30594
440923d2
700c50ad
c2d240a6
323c4086
700f231b
0286275c
0108931c
975c06b4
80060066
04b3c026
0108101c
393c3cce
43c3ef80
fef34364
686c2bc3
001c6ccc
011c0bb4
20260000
353c3664
073c0010
24c33f9d
01ff431c
201c0335
23640200
180c353c
4cce7d80
43c37120
c0254364
536456c3
e1948007
0296675c
31c33c2b
1d806205
28c31c4f
2c544007
24c37ccb
26143ae4
45d22cc3
2ac31cc3
08cbb0bc
3c4c3ac3
18c30c80
23c37ccb
b0bc2aa4
3ccb08cb
3aa431c3
40268384
423c0233
323c0010
bd80180c
4e1d073c
253c18c3
b0bc063e
540b08cb
24c38284
26e42364
2006ef14
07c33c2f
f8760196
08040f56
0736f016
80c3fd96
02c3a1c3
13c30364
e0061364
34c347c3
68f237a3
a8cb28c3
7e0535c3
236423c3
373c0113
6e000067
58c360c5
359d253c
053402e4
901c61c3
0af30000
03c36120
80270364
80260354
373c00f3
60b70010
00417f5c
00078006
fdb3db94
37a334c3
58c36cf2
6280b48c
0100133c
a8cb28c3
7e0535c3
02336c20
0037373c
60856e00
223c28c3
21003a1d
0067373c
60c56e00
553c58c3
7420359d
236423c3
236402c3
023526e4
50c306c3
0ac35364
25c30984
08cbb0bc
033465e4
0093c006
63c37aa0
80276364
273c0894
40770010
00217f5c
00d38006
0010243c
4f5c4037
29c30001
93c37500
00069364
b994c007
e0760396
08040f56
3f36f016
2177fa96
c364c3c3
02231f5c
02413f5c
0cc36137
83c36800
00048364
600738c3
000af2dc
1110301c
0000311c
6c0c25d2
00a66e8c
6c0c0093
00866e8c
00812f5c
366412c3
000760c3
0009b2dc
408cd0c3
620f6006
0100383c
680c638e
601b383c
901c680f
b9c30000
79c3a9c3
00f0301c
33643ca4
09c36037
27940007
831c8017
05b400f0
3ca438c3
436443c3
388c0cc3
033c6080
41570100
1b8412c3
b0bc24c3
0cc308cb
23c37000
38cb2364
620531c3
78ce6980
612008c3
836483c3
0010373c
7f5c60f7
0a330061
1110001c
0000011c
6c4c600c
401c6c6c
411c0bb4
6ccc0000
200604c3
50c33664
301c0ff2
311c0ef0
6c0c0000
163c100c
36640040
62bc0f86
d5c30a77
3a3c07f3
6f800037
063c6085
28c33b9d
336438c3
0200331c
201c0335
42c30200
05c34364
12c34157
24c31b84
08cbb0bc
00673a3c
60c56f80
371d463c
622008c3
836483c3
0a94e027
00100a3c
1f5c00b7
a1c30041
e006a264
373c00d3
60770010
00217f5c
0cd208c3
70801bc3
b364b3c3
0010393c
936493c3
d01cefb3
0dc30000
fc760696
08040f56
0f36f016
70c3fd96
826481c3
8100402b
706c2050
242b333c
301c706f
311c1110
4c0c0000
48d0a80c
0bb4301c
0000311c
700c6ed0
f000341c
5000331c
001c0454
2193009b
200675ec
1000111c
64d23183
20066b4c
29c33664
610768cb
331c0c54
09540608
dd86101c
0000111c
32e421c3
000f74dc
0a0502bc
570b60c3
0056323c
7f327fe5
18c36cd2
f8bc2ad2
60c30a04
01a1255c
801c40b7
03930003
11546007
6ff238c3
0229155c
11542007
00478f5c
01a1255c
602643f2
801c60b7
01530000
20b72006
831c82c3
04540003
60b76006
09c383c3
40c616c3
08cbeabc
0060393c
52940007
16c303c3
eabc40c6
000708cb
000b72dc
25291ac3
19542007
0bb4301c
0000311c
6e0c6c2c
12c34dc9
323c4de9
6df240ac
65891ac3
04946047
658c1bc3
2bc33664
1ac369ac
366404ab
133c75ec
20770014
3b942007
400653c3
0004211c
a0075283
3f5c7354
704d0021
0003831c
501c5f94
511c1110
740c0000
04a4335c
2f5c07c3
12c30041
30c33664
60073264
60264f54
740c704d
0484335c
17c30057
00573664
03c30e73
40c616c3
08cbeabc
5a540007
440919c3
341c32c3
60070001
75ec5854
0014233c
4cd24037
1110301c
0000311c
335c6c0c
00060484
366417c3
53c30673
111c2006
51830004
2e54a007
00012f5c
831c504d
1a940003
1110501c
0000511c
335c740c
07c304a4
00412f5c
366412c3
326430c3
60266bd2
740c704d
0484335c
17c30017
00173664
301c05f3
311c1110
6c0c0000
04c4335c
2f5c07c3
12c30041
00063664
301c0433
311c1110
6c0c0000
04c4335c
2f5c07c3
12c30041
05c33664
706c0273
323c4026
706f241b
7ccb0026
001c6bf2
62bc00b3
706c0a77
323c4026
706f241b
039602c3
0f56f076
00000804
00f34006
0014303c
488062d2
21120132
02c31af2
00000804
40c33016
602601c3
41120073
20e46112
6bd20c34
fa154007
02e40113
01200314
613213a3
00534132
78f22006
01c382f2
08040c56
50c37016
62c341c3
0b0d113c
0b0d223c
0a7bc0bc
8007a4d2
01330b15
800725c3
40260215
f88c363c
025423e4
0e5600c4
00000804
50c33016
436441c3
20262364
323c0133
23c3080c
313c2364
13c3080c
24e41364
2fd21034
316432c3
f2156007
42e40153
71200514
436443c3
213201a3
00534132
36f20006
04c3a2d2
08040c56
50c37016
416441c3
616462c3
0b0d143c
0b0d263c
0a7bf4bc
a4d20364
0b158007
25c30133
02158007
363c4026
23e4f88c
00c40254
08040e56
316430c3
216421c3
13c30006
0a7c1abc
00000804
336430c3
236421c3
13c30006
0a7bf4bc
00000804
316430c3
216421c3
13c30026
0a7c1abc
00000804
21c330c3
13c30026
0a7bf4bc
00000804
203c3016
313c0b0d
141d0b0d
513c4230
bf32001c
0354a007
005304c4
0c5604c3
00000804
203c1016
313c0b0d
341d0b0d
1f324230
03540007
005304c4
085604c3
00000804
40c31016
111c2006
c2bc4700
00070a98
04c30f74
111c2006
08bc4700
04bc0a95
301c0a94
311c8000
01800000
04c30093
0a9404bc
08040856
11c4fc96
0b0d303c
7f3233c4
25a000c4
08040496
fc961016
400741c3
64061654
20072d20
600607d4
31c46077
308d343c
343c0133
6077208d
100d343c
208d203c
603732a3
80570017
049614c3
08040856
fc961016
400740c3
64061654
00070d20
600607d4
30c46037
300d343c
343c0133
6037200d
008d343c
200d213c
607732a3
20578017
049604c3
08040856
fc961016
400741c3
64061754
20072d20
343c08d4
6077f90c
343c31c4
0133310d
210d343c
343c6077
203c100d
32a3208d
00176037
14c38057
08560496
00000804
4406fe96
01c323d2
60064006
0b8d303c
02960d00
00000804
fc961016
13e440c3
13e40974
42e409d4
00260514
053542e4
00060073
00460053
08560496
00000804
fc961016
13e440c3
13e40914
42e409b4
00260514
053542e4
00060073
00460053
08560496
00000804
3f36f016
c0c3fc96
b2c351c3
df5c73c3
32c301e4
62f237a3
75e40013
75e405b4
b0e40c94
1dc30a35
25d26dc3
88112dc3
c006a82f
0ad386c3
c4063cc3
35c3a3d2
8006c006
233c24c3
1bc30b8d
e3d20406
04c317c3
34c38006
0b8d313c
61805900
92a493c3
15c30cc3
a4bc29c3
64c30a7c
363c84c3
483cf88c
c11209ac
71e484c3
71e417b4
b0e40394
263c13b4
60260010
021426e4
62c36006
848483c3
81a03bc3
40e44026
400602b4
04c367a0
29c32d20
14544007
ffff921c
f88c303c
09aca13c
080c403c
15c30cc3
a4bc29c3
303c0a7c
04c30014
1ac303a3
3dc3f9b3
0c0f63d2
06c32c2f
049618c3
0f56fc76
70160804
41c3fb96
00f763c3
40772137
a00660b7
0a1545e4
202600c4
10c302f2
6ca034c4
613700f7
6097bfe6
0a156007
22c455e3
42f22026
36c412c3
40776ca0
600660b7
00d76037
40572117
34bc6097
20c30a7d
a7d231c3
202602c4
10c302f2
2ca033c4
0e560596
00000804
ff961016
80378006
0a7d34bc
08560196
00000804
f9967016
53c341c3
21b70177
613740f7
46e4c006
00c40a15
02f22026
34c410c3
01776ca0
dfe661b7
60076117
22c40915
42f22026
35c412c3
40f76ca0
3f3c6137
60370040
21970157
611740d7
0a7d34bc
0097cbd2
23c46057
42f22026
30c412c3
40776ca0
005760b7
07962097
08040e56
fd961016
00404f3c
34bc8037
00570a7d
03962097
08040856
0136f016
50c3fe96
803c41c3
713c808c
21c3808c
023c2364
35c3828d
133c3364
333c728d
233c228d
30c3808c
ffff341c
203ccd00
313c808c
4980808c
828d373c
141c4980
7880ffff
043c7032
2980528d
80760296
08040f56
fa96f016
52c370c3
43c361c3
2ebc12c3
273c0a7e
353c428d
6980628d
06962580
08040f56
13bc301c
0000311c
4c0f4006
6c4f4c2f
301c6c6f
311c13b0
4c0f0000
13ac301c
0000311c
301c4c0f
311c13b4
4c0f0000
13b8301c
0000311c
08044c0f
0336f016
0e2440c3
f52480c3
10fc301c
0000311c
343c4c0c
6e20f90c
033c496c
2664f88c
02b480e7
343c8106
5f860030
533c3283
301c0080
311c13bc
4c4c0000
282c0233
0d7415e4
13bc601c
0000611c
39e496c3
0c2c0554
14e440c3
32c30215
601c484c
611c13bc
96c30000
ea9429e4
111343c3
25e4502c
000843dc
101c6aa0
111c10fc
62070000
d1803135
240cfa80
7c0c0006
029432e4
656c0026
702c3664
702f6ea0
35c4780f
0006782f
301c1c0f
311c13ac
2c0c0000
8c0f9480
13b0201c
0000211c
34e4680c
880f0215
13b4201c
0000211c
6025680c
063c680f
383c0080
60074004
f3245d54
b1000b73
0006240c
32e4740c
00260294
3664656c
10fc301c
0000311c
00064c0c
6c4c706c
029434e4
696c0026
301c3664
311c10fc
4c0c0000
704c0006
34e46c6c
00260294
3664696c
704c506c
704c684f
201c4c6f
211c13ac
702c0000
2f00c80c
201c280f
211c13b4
680c0000
680f6025
13b0201c
0000211c
31e4680c
280f0215
33c4702c
0006702f
383c140f
62d24004
043cf324
02130080
101c904c
111c13bc
21c30000
34dc42e4
383cfff7
03c34004
f32463d2
c0760006
08040f56
60c3f016
f524ee24
ff80503c
13b8201c
0000211c
6025680c
401c680f
411c10fc
500c0000
0b0d303c
496c33c4
f88c033c
900c2664
742c0006
021530e4
716c0026
301c3664
311c10fc
4c0c0000
742c0006
758133c4
002662f2
3664696c
13ac201c
0000211c
880c742c
280f2e00
10fc401c
0000411c
21e3700c
023c6d6c
3664f88c
0007140c
d42c1154
4006300c
6c2c7420
029430e4
656c4026
366402c3
b420140c
6f20742c
500c0673
13bc301c
0000311c
6c4c6c6c
13bc101c
0000111c
34e441c3
00260294
3664696c
10fc301c
0000311c
00064c0c
13bc301c
0000311c
6c6c6c4c
13bc101c
0000111c
34e441c3
00260294
3664696c
13bc301c
0000311c
4c6c780f
ac6f546f
742ca84f
742f33c4
9700d42c
4007502c
301c31f4
311c10fc
2c0c0000
71010006
029432e4
656c0026
301c3664
311c10fc
4c0c0000
706c0006
34e46c4c
00260294
3664696c
